* NGSPICE file created from team_08.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

.subckt team_08 clk en gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3]
+ gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0]
+ gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16]
+ gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22]
+ gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29]
+ gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XFILLER_0_20_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4654__B allocation.game.controller.drawBlock.y_start\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_7963_ allocation.game.controller.v\[2\] allocation.game.controller.v\[1\] allocation.game.controller.v\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3476_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6914_ _2683_ _2684_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__nor2_1
X_7894_ _3427_ vssd1 vssd1 vccd1 vccd1 _3428_ sky130_fd_sc_hd__inv_2
X_6845_ allocation.game.cactus2size.clock_div_inst0.counter\[11\] allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ _2634_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7590__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6776_ allocation.game.cactus2size.clock_div_inst1.counter\[1\] allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ _2592_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__o21ai_1
X_9495_ clknet_leaf_12_clk _0395_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.internalSck
+ sky130_fd_sc_hd__dfxtp_1
X_5727_ _1649_ _1650_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__xnor2_1
X_8515_ net51 net48 _3328_ _3966_ _3346_ vssd1 vssd1 vccd1 vccd1 _3967_ sky130_fd_sc_hd__a41o_1
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8446_ _3289_ _3324_ vssd1 vssd1 vccd1 vccd1 _3899_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5658_ _0761_ _0887_ _1538_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__and3_1
X_4609_ net262 net231 _0511_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__a21o_1
X_8377_ allocation.game.dinoJump.next_dinoY\[0\] _0530_ _0534_ _0538_ vssd1 vssd1
+ vccd1 vccd1 _3838_ sky130_fd_sc_hd__and4_1
X_5589_ _1509_ _1512_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7328_ net223 net151 _0616_ _2313_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7259_ allocation.game.controller.init_module.delay_counter\[0\] _2926_ vssd1 vssd1
+ vccd1 vccd1 _2929_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout75_A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9432__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8373__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8052__A _4459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4960_ _0705_ _0706_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4891_ _0725_ _0814_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6630_ _2496_ net150 _2495_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[20\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_27_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6561_ _2448_ _2449_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[19\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8300_ net81 _2253_ vssd1 vssd1 vccd1 vccd1 _3766_ sky130_fd_sc_hd__nor2_1
X_5512_ _1426_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__nor2_1
X_6492_ _0417_ allocation.game.controller.drawBlock.state\[0\] allocation.game.controller.drawBlock.state\[3\]
+ _0606_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a22o_1
XANTENNA__9305__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9280_ clknet_leaf_0_clk _0095_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8231_ allocation.game.lcdOutput.tft.remainingDelayTicks\[7\] _2987_ vssd1 vssd1
+ vccd1 vccd1 _3714_ sky130_fd_sc_hd__xor2_1
X_5443_ _1341_ _1363_ _1365_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__and3_1
X_8162_ allocation.game.controller.state\[2\] _3658_ _0627_ vssd1 vssd1 vccd1 vccd1
+ _3659_ sky130_fd_sc_hd__o21a_1
X_5374_ _1202_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nand2_1
X_7113_ _2757_ _2824_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout138 _3461_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_1
X_8093_ net242 net281 _2413_ vssd1 vssd1 vccd1 vccd1 _3597_ sky130_fd_sc_hd__or3_4
Xfanout105 _0672_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_1
Xfanout127 allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1 vccd1
+ net127 sky130_fd_sc_hd__buf_1
XFILLER_0_11_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout116 _3182_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_2
X_7044_ allocation.game.controller.drawBlock.idx\[2\] _0443_ allocation.game.controller.drawBlock.idx\[1\]
+ allocation.game.controller.drawBlock.idx\[4\] vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__a31o_1
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_2
X_8995_ net142 net59 _4099_ _4107_ _4108_ vssd1 vssd1 vccd1 vccd1 _4444_ sky130_fd_sc_hd__a2111o_1
X_7946_ net231 allocation.game.controller.v\[5\] allocation.game.controller.v\[4\]
+ allocation.game.controller.v\[7\] vssd1 vssd1 vccd1 vccd1 _3460_ sky130_fd_sc_hd__or4_2
XFILLER_0_49_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7695__B net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7877_ _3415_ vssd1 vssd1 vccd1 vccd1 _3416_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6828_ allocation.game.cactus2size.clock_div_inst0.counter\[5\] _2625_ vssd1 vssd1
+ vccd1 vccd1 _2627_ sky130_fd_sc_hd__and2_1
XANTENNA__5496__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6759_ allocation.game.cactus1size.clock_div_inst0.counter\[10\] _2578_ _2580_ vssd1
+ vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9478_ clknet_leaf_7_clk _0385_ net187 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.v\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8429_ _3881_ vssd1 vssd1 vccd1 vccd1 _3882_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout78_X net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8830__A3 _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4575__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5801__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9328__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8510__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9478__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6030__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7560__S net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8282__B2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8282__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5090_ _0731_ _0949_ _0995_ _0997_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__a31o_1
X_5992_ _1913_ _1914_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__xnor2_1
X_8780_ _3486_ _3760_ vssd1 vssd1 vccd1 vccd1 _4230_ sky130_fd_sc_hd__nand2_1
X_7800_ _2861_ _3355_ vssd1 vssd1 vccd1 vccd1 _3362_ sky130_fd_sc_hd__or2_2
X_4943_ _0866_ _0867_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__nor2_1
X_7731_ _3248_ net46 vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__and2_2
XFILLER_0_8_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7662_ allocation.game.lcdOutput.framebufferIndex\[8\] _3213_ net56 _3210_ vssd1
+ vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4874_ _0543_ _0572_ _0768_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__nand3_2
X_6613_ allocation.game.cactusMove.count\[13\] allocation.game.cactusMove.count\[14\]
+ _2482_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__and3_1
X_9401_ clknet_leaf_17_clk _0311_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7593_ net144 _3169_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9332_ clknet_leaf_6_clk _0115_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_6544_ _2437_ _2438_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[13\]
+ sky130_fd_sc_hd__nor2_1
X_6475_ allocation.game.scoreCounter.clock_div.counter\[13\] allocation.game.scoreCounter.clock_div.counter\[10\]
+ allocation.game.scoreCounter.clock_div.counter\[14\] vssd1 vssd1 vccd1 vccd1 _2390_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9263_ clknet_leaf_2_clk _0055_ net189 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_8214_ _0624_ _3702_ net113 vssd1 vssd1 vccd1 vccd1 _3703_ sky130_fd_sc_hd__a21oi_1
X_5426_ _1202_ _1298_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__or2_1
X_9194_ clknet_leaf_12_clk net362 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.cs
+ sky130_fd_sc_hd__dfxtp_1
X_8145_ _0612_ _2524_ vssd1 vssd1 vccd1 vccd1 _3644_ sky130_fd_sc_hd__nand2_1
X_5357_ _1280_ _1281_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__nor2_1
X_8076_ net140 _3579_ _3581_ _3582_ vssd1 vssd1 vccd1 vccd1 _3583_ sky130_fd_sc_hd__o22a_1
XANTENNA__8273__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5288_ _1195_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7027_ _0439_ allocation.game.scoreCounter.bcd_tens\[2\] _2749_ vssd1 vssd1 vccd1
+ vccd1 _2754_ sky130_fd_sc_hd__o21a_1
X_8978_ _0678_ net98 net76 _0651_ _4426_ vssd1 vssd1 vccd1 vccd1 _4427_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_2_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7929_ _3452_ vssd1 vssd1 vccd1 vccd1 _3453_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8984__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7380__S _2973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5078__A1 _0938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4825__A1 _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9150__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7555__S net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4590_ _0523_ _0524_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4646__A_N allocation.game.controller.drawBlock.y_start\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6260_ _1983_ _2107_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5211_ _0846_ _1078_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__nor2_1
X_6191_ _2114_ _2115_ _1763_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5142_ _1065_ _1066_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5073_ _0985_ _0996_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__xnor2_1
X_8901_ _4350_ _3916_ _4333_ vssd1 vssd1 vccd1 vccd1 _4351_ sky130_fd_sc_hd__or3b_1
XANTENNA__8415__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8832_ net38 _4279_ _4281_ net36 vssd1 vssd1 vccd1 vccd1 _4282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4662__B allocation.game.controller.drawBlock.y_end\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5975_ _1790_ _1793_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__nand2_1
X_8763_ net268 _4212_ vssd1 vssd1 vccd1 vccd1 _4213_ sky130_fd_sc_hd__nand2_1
X_4926_ _0840_ _0845_ _0849_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_47_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7714_ net39 net41 vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__nand2_1
X_8694_ _4137_ _4139_ _4142_ _4144_ vssd1 vssd1 vccd1 vccd1 _4145_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4857_ _0763_ _0781_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7645_ _3194_ _3195_ _3206_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7576_ allocation.game.cactus1size.lfsr1\[1\] allocation.game.cactus1size.lfsr1\[0\]
+ allocation.game.cactus1size.clock_div_inst0.clk1 vssd1 vssd1 vccd1 vccd1 _3160_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9315_ clknet_leaf_6_clk _0122_ net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4788_ _0563_ _0711_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__or2_1
X_6527_ net393 _2425_ _2427_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[7\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6458_ net222 _2311_ _2374_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9246_ clknet_leaf_1_clk net395 net176 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6389_ _0415_ net218 vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__and2_1
X_5409_ _0751_ _0949_ _1333_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_8_Left_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9177_ clknet_leaf_18_clk _0239_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.initSeqCounter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_8128_ net112 _0689_ vssd1 vssd1 vccd1 vccd1 _3628_ sky130_fd_sc_hd__nor2_1
XANTENNA__7988__X _3500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8059_ _0509_ _3565_ vssd1 vssd1 vccd1 vccd1 _3567_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4807__A1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5760_ _0769_ _0905_ _0907_ _0777_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__a22o_1
XANTENNA__8960__A2 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4711_ net226 allocation.game.cactusMove.x_dist\[4\] _0637_ vssd1 vssd1 vccd1 vccd1
+ _0638_ sky130_fd_sc_hd__a21oi_2
X_5691_ _1613_ _1614_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4642_ _0545_ _0571_ _0544_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__a21o_2
XANTENNA__8173__B1 _3609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7430_ _3046_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4573_ _0507_ _0508_ _0509_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9046__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7361_ allocation.game.lcdOutput.tft.remainingDelayTicks\[22\] allocation.game.lcdOutput.tft.remainingDelayTicks\[23\]
+ _2998_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__or3_2
X_7292_ net474 _2947_ _2950_ _2928_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__o211a_1
X_6312_ allocation.game.controller.drawBlock.state\[2\] _0606_ _2234_ _2236_ vssd1
+ vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9100_ clknet_leaf_9_clk _0196_ net198 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight1\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9031_ clknet_leaf_4_clk _0156_ net185 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6243_ _2119_ _2120_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4657__B allocation.game.controller.drawBlock.y_end\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6174_ _2078_ _2097_ _2066_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__a21o_1
X_5125_ _0797_ _1049_ _1013_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout192_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5056_ _0979_ _0976_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_28_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8400__A1 allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8815_ _4253_ _4254_ _4263_ _4264_ vssd1 vssd1 vccd1 vccd1 _4265_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8746_ net227 net257 net164 net142 vssd1 vssd1 vccd1 vccd1 _4197_ sky130_fd_sc_hd__a31oi_2
X_5958_ _1879_ _1880_ _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__nand3_1
X_4909_ _0794_ _0804_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__nand2_4
XFILLER_0_30_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5889_ _0723_ net86 vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__nor2_1
X_8677_ net120 _4127_ vssd1 vssd1 vccd1 vccd1 _4128_ sky130_fd_sc_hd__nor2_1
XANTENNA__5517__A2 _0886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7628_ _3178_ _3179_ _3183_ _3189_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__o31a_1
X_7559_ net327 allocation.game.lcdOutput.tft.spi.data\[6\] net256 vssd1 vssd1 vccd1
+ vccd1 _0247_ sky130_fd_sc_hd__mux2_1
X_9229_ clknet_leaf_22_clk _0026_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold30 allocation.game.lcdOutput.tft.spi.tft_dc vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 allocation.game.lcdOutput.tft.spi.data\[1\] vssd1 vssd1 vccd1 vccd1 net364
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 allocation.game.scoreCounter.clock_div.counter\[24\] vssd1 vssd1 vccd1 vccd1
+ net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold52 allocation.game.lcdOutput.tft.remainingDelayTicks\[17\] vssd1 vssd1 vccd1
+ vccd1 net375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 allocation.game.dinoJump.dinoDelay\[17\] vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4583__A _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold85 allocation.game.controller.drawBlock.x_end\[5\] vssd1 vssd1 vccd1 vccd1 net408
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 allocation.game.dinoJump.count\[6\] vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6650__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5205__A1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9069__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7902__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4758__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6930_ net160 _2693_ _2694_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__nor3_1
XFILLER_0_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6861_ allocation.game.cactusDist.clock_div_inst1.counter\[1\] allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ allocation.game.cactusDist.clock_div_inst1.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2649_ sky130_fd_sc_hd__nand3_1
X_5812_ net71 _0903_ _1684_ _1685_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__a22o_1
X_8600_ net46 _4044_ _4045_ _4050_ _4049_ vssd1 vssd1 vccd1 vccd1 _4051_ sky130_fd_sc_hd__o41a_1
X_6792_ allocation.game.cactus2size.clock_div_inst1.counter\[7\] _2601_ net158 vssd1
+ vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5743_ _1627_ _1628_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8531_ _3915_ _3970_ _3981_ _3967_ _3982_ vssd1 vssd1 vccd1 vccd1 _3983_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8146__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5674_ _1597_ _1598_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__nand2_1
X_8462_ net114 _3914_ vssd1 vssd1 vccd1 vccd1 _3915_ sky130_fd_sc_hd__nor2_1
X_8393_ _3841_ _3850_ _3848_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a21oi_1
X_4625_ _0553_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__nand2b_1
X_7413_ allocation.game.lcdOutput.tft.state\[0\] net55 _3030_ _3033_ vssd1 vssd1 vccd1
+ vccd1 _3034_ sky130_fd_sc_hd__and4_1
X_4556_ _4457_ allocation.game.controller.v\[1\] vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7344_ allocation.game.lcdOutput.tft.remainingDelayTicks\[2\] _2983_ vssd1 vssd1
+ vccd1 vccd1 _2984_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout205_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4487_ allocation.game.controller.init_module.delay_counter\[23\] vssd1 vssd1 vccd1
+ vccd1 _0427_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7275_ net477 _2937_ _2939_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_38_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6226_ _2147_ _2150_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__xnor2_1
X_9014_ net255 vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7672__A2 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6157_ net110 _0894_ _2081_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout195_X net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8082__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5108_ _1026_ _1031_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6632__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6088_ _1972_ _1984_ _2008_ _2012_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__a31o_1
X_5039_ _0880_ _0882_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__a21oi_1
X_9527__321 vssd1 vssd1 vccd1 vccd1 net321 _9527__321/LO sky130_fd_sc_hd__conb_1
XFILLER_0_36_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7219__A _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8729_ net121 _4179_ vssd1 vssd1 vccd1 vccd1 _4180_ sky130_fd_sc_hd__nor2_1
XANTENNA__9361__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput7 net7 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__clkbuf_4
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5390_ _1312_ _1314_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4488__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7060_ allocation.game.controller.drawBlock.x_end\[0\] _2777_ _2779_ allocation.game.controller.drawBlock.y_end\[0\]
+ _2776_ vssd1 vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__a221o_1
X_6011_ _1893_ _1894_ _1886_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9234__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7962_ _3470_ _3471_ _3472_ _3474_ vssd1 vssd1 vccd1 vccd1 _3475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6913_ allocation.game.cactusDist.clock_div_inst0.counter\[5\] _2681_ net155 vssd1
+ vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__o21ai_1
X_7893_ allocation.game.controller.drawBlock.counter\[7\] allocation.game.controller.drawBlock.counter\[8\]
+ _3423_ vssd1 vssd1 vccd1 vccd1 _3427_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9384__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout155_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6844_ allocation.game.cactus2size.clock_div_inst0.counter\[10\] _2634_ allocation.game.cactus2size.clock_div_inst0.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__a21oi_1
X_6775_ allocation.game.cactus2size.clock_div_inst1.counter\[0\] _2592_ vssd1 vssd1
+ vccd1 vccd1 _0062_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5726_ _1650_ _1649_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__nand2b_1
X_8514_ _3289_ _3303_ vssd1 vssd1 vccd1 vccd1 _3966_ sky130_fd_sc_hd__nor2_1
X_9494_ clknet_leaf_16_clk _0394_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.r_floor
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8445_ _3303_ _3366_ _3893_ _3365_ net96 vssd1 vssd1 vccd1 vccd1 _3898_ sky130_fd_sc_hd__o32a_1
X_5657_ _0761_ _0887_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout110_X net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8376_ allocation.game.controller.v\[0\] net84 vssd1 vssd1 vccd1 vccd1 _3837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4608_ net260 _0481_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__or2_1
X_5588_ _1509_ _1512_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__or2_1
X_4539_ allocation.game.dinoJump.count\[6\] allocation.game.dinoJump.count\[8\] allocation.game.dinoJump.count\[10\]
+ allocation.game.dinoJump.count\[7\] vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__or4b_1
X_7327_ _0616_ _2972_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__nand2_4
X_7258_ _2821_ _2926_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__nand2_1
X_6209_ _1118_ _2133_ _1117_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7189_ _0472_ _2873_ _2875_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout68_A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5022__A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6081__B2 _0729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6788__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9107__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9257__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4890_ _0725_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6560_ net471 _2447_ net90 vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5511_ _0710_ _0717_ _0718_ _1435_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6491_ _2235_ _2234_ net412 _0417_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__a2bb2o_1
X_8230_ _3025_ _3032_ _3713_ _3001_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__a22o_1
X_5442_ _1336_ _1358_ _1360_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__a21o_1
X_8161_ allocation.game.controller.state\[7\] _3465_ vssd1 vssd1 vccd1 vccd1 _3658_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5373_ _0975_ _1201_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7112_ _2820_ _2823_ allocation.game.controller.init_module.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _2824_ sky130_fd_sc_hd__o21ai_1
X_8092_ net230 net203 vssd1 vssd1 vccd1 vccd1 _3596_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_35_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7043_ _2762_ _2763_ allocation.game.controller.drawBlock.idx\[3\] _0444_ vssd1 vssd1
+ vccd1 vccd1 _2764_ sky130_fd_sc_hd__o2bb2a_1
Xfanout106 _0480_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout117 net119 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout128 allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1 vccd1
+ net128 sky130_fd_sc_hd__buf_2
Xfanout139 _3461_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_8994_ net142 net59 net52 _0655_ _4442_ vssd1 vssd1 vccd1 vccd1 _4443_ sky130_fd_sc_hd__o221a_1
X_7945_ net370 _0695_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7876_ allocation.game.controller.drawBlock.counter\[0\] allocation.game.controller.drawBlock.counter\[1\]
+ allocation.game.controller.drawBlock.counter\[2\] allocation.game.controller.drawBlock.counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _3415_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6827_ _2625_ _2626_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6758_ allocation.game.cactus1size.clock_div_inst0.counter\[10\] _2578_ net160 vssd1
+ vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_21_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9477_ clknet_leaf_7_clk _0384_ net194 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.v\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_6689_ _2534_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__inv_2
X_5709_ _1619_ _1632_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8428_ _3303_ _3370_ vssd1 vssd1 vccd1 vccd1 _3881_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8359_ _3814_ _3821_ allocation.game.controller.drawBlock.y_end\[6\] net201 vssd1
+ vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold160 allocation.game.controller.init_module.delay_counter\[7\] vssd1 vssd1 vccd1
+ vccd1 net483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8028__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8579__B1 _3996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9505__290 vssd1 vssd1 vccd1 vccd1 _9505__290/HI net290 sky130_fd_sc_hd__conb_1
XFILLER_0_3_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6030__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4766__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5991_ net87 _0900_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4942_ _0833_ _0865_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__and2_1
X_7730_ _3237_ _3249_ vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7661_ allocation.game.lcdOutput.framebufferIndex\[7\] _3213_ _3222_ vssd1 vssd1
+ vccd1 vccd1 _3223_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6612_ allocation.game.cactusMove.count\[12\] allocation.game.cactusMove.count\[13\]
+ _2480_ allocation.game.cactusMove.count\[14\] vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__a31o_1
X_4873_ _0710_ net79 vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__or2_4
X_9400_ clknet_leaf_17_clk _0310_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7592_ allocation.game.cactus2size.lfsr2\[1\] allocation.game.cactus2size.lfsr2\[0\]
+ allocation.game.cactus2size.clock_div_inst1.clk1 vssd1 vssd1 vccd1 vccd1 _3169_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9422__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9331_ clknet_leaf_6_clk _0114_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_6543_ allocation.game.dinoJump.dinoDelay\[13\] _2436_ net90 vssd1 vssd1 vccd1 vccd1
+ _2438_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6474_ allocation.game.scoreCounter.clock_div.counter\[18\] allocation.game.scoreCounter.clock_div.counter\[17\]
+ _2387_ _2388_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9262_ clknet_leaf_2_clk _0054_ net191 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_8213_ net219 _0623_ net218 vssd1 vssd1 vccd1 vccd1 _3702_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout118_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5425_ _1349_ _1347_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__nand2b_1
X_9193_ clknet_leaf_15_clk _0254_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.tft_sdi
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8144_ _0415_ _3634_ vssd1 vssd1 vccd1 vccd1 _3643_ sky130_fd_sc_hd__nand2_1
X_5356_ _1274_ _1277_ _1279_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8075_ _0541_ _3565_ _3580_ net136 vssd1 vssd1 vccd1 vccd1 _3582_ sky130_fd_sc_hd__a31o_1
X_5287_ _1208_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__xnor2_1
X_7026_ allocation.game.scoreCounter.bcd_tens\[1\] allocation.game.scoreCounter.bcd_tens\[0\]
+ _2753_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__or3_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8977_ net120 _3647_ _3190_ _0679_ vssd1 vssd1 vccd1 vccd1 _4426_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7928_ allocation.game.controller.drawBlock.counter\[17\] allocation.game.controller.drawBlock.counter\[18\]
+ _3447_ vssd1 vssd1 vccd1 vccd1 _3452_ sky130_fd_sc_hd__and3_1
XANTENNA__5300__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7859_ allocation.game.controller.drawBlock.idx\[1\] _3402_ _3403_ _3404_ vssd1 vssd1
+ vccd1 vccd1 _0296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9529_ net323 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6131__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4586__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4825__A2 _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4873__X _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9445__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5210_ _1132_ _1134_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5710__B1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6190_ _1761_ _1762_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__xnor2_1
X_5141_ _0754_ _0772_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__xnor2_1
X_5072_ _0985_ _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8900_ _4347_ _4349_ vssd1 vssd1 vccd1 vccd1 _4350_ sky130_fd_sc_hd__nor2_1
X_8831_ _0468_ _4277_ _4280_ vssd1 vssd1 vccd1 vccd1 _4281_ sky130_fd_sc_hd__o21ai_1
X_8762_ _4458_ _3486_ vssd1 vssd1 vccd1 vccd1 _4212_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7713_ _3258_ _3273_ vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__or2_1
X_5974_ _1790_ _1793_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ _0840_ _0845_ _0849_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_47_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8693_ _4132_ _4133_ _4143_ _4129_ _4128_ vssd1 vssd1 vccd1 vccd1 _4144_ sky130_fd_sc_hd__a311o_1
X_4856_ net103 _0740_ _0743_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__mux2_2
X_7644_ _3185_ _3186_ _3202_ _3184_ vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7575_ allocation.game.cactus1size.lfsr1\[0\] _3158_ _3159_ vssd1 vssd1 vccd1 vccd1
+ _0257_ sky130_fd_sc_hd__o21ai_1
X_9314_ clknet_leaf_5_clk net382 net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4787_ _0563_ _0711_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6526_ allocation.game.dinoJump.dinoDelay\[7\] _2425_ _2415_ vssd1 vssd1 vccd1 vccd1
+ _2427_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6457_ net222 _2311_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5790__A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9245_ clknet_leaf_1_clk _0062_ net177 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6388_ net222 _2311_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__nor2_1
X_5408_ _1331_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9176_ clknet_leaf_16_clk _0238_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.initSeqCounter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8127_ _0651_ _3614_ _3626_ _0419_ vssd1 vssd1 vccd1 vccd1 _3627_ sky130_fd_sc_hd__a211oi_1
X_5339_ _1253_ _1256_ _1262_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__nand3_1
XANTENNA__9318__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8058_ _3563_ _3564_ net139 vssd1 vssd1 vccd1 vccd1 _3566_ sky130_fd_sc_hd__a21o_1
XANTENNA__4807__A2 _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7009_ _0450_ _0451_ _2736_ _2743_ vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__a31oi_1
XANTENNA__8606__A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout50_A _3228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9468__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4747__C net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7566__S _2526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4710_ _0635_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__and2b_1
X_5690_ _1614_ _1613_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4641_ _0548_ _0570_ _0547_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4572_ _0507_ _0508_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__and3_1
X_7360_ allocation.game.lcdOutput.tft.remainingDelayTicks\[23\] _2999_ vssd1 vssd1
+ vccd1 vccd1 _3000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7291_ _2949_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__inv_2
X_6311_ net236 allocation.game.controller.drawBlock.state\[3\] _0606_ vssd1 vssd1
+ vccd1 vccd1 _2236_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9030_ clknet_leaf_4_clk _0155_ net187 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6242_ _1531_ _2121_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6173_ _2078_ _2097_ _2066_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__a21oi_1
X_5124_ _1045_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout185_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5055_ _0976_ _0979_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__and2b_1
XANTENNA__4673__B allocation.game.controller.drawBlock.y_start\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8814_ net44 _4261_ vssd1 vssd1 vccd1 vccd1 _4264_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4960__Y _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5957_ _1820_ _1881_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__xnor2_1
X_8745_ net227 _0654_ _3594_ vssd1 vssd1 vccd1 vccd1 _4196_ sky130_fd_sc_hd__mux2_1
X_4908_ _0778_ _0832_ _0798_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__mux2_2
XFILLER_0_30_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8676_ _0675_ _4122_ _4126_ vssd1 vssd1 vccd1 vccd1 _4127_ sky130_fd_sc_hd__o21ai_1
X_5888_ net141 _0888_ _1768_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__or3b_1
X_7627_ _2843_ _3180_ _3188_ vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_44_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4839_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7558_ net346 net345 allocation.game.lcdOutput.tft.spiDataSet vssd1 vssd1 vccd1 vccd1
+ _0246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7489_ net247 _3102_ vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__nor2_1
X_6509_ allocation.game.dinoJump.dinoDelay\[1\] allocation.game.dinoJump.dinoDelay\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__nand2_1
X_9228_ clknet_leaf_21_clk _0025_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5025__A _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9159_ clknet_leaf_18_clk _0221_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold31 _0253_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold20 allocation.game.lcdOutput.tft.spi.data\[2\] vssd1 vssd1 vccd1 vccd1 net343
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold42 allocation.game.lcdOutput.tft.remainingDelayTicks\[2\] vssd1 vssd1 vccd1 vccd1
+ net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 allocation.game.dinoJump.dinoDelay\[11\] vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 allocation.game.lcdOutput.tft.remainingDelayTicks\[19\] vssd1 vssd1 vccd1
+ vccd1 net376 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9290__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold97 allocation.game.controller.init_module.delay_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 allocation.game.controller.drawBlock.y_start\[1\] vssd1 vssd1 vccd1 vccd1
+ net409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 allocation.game.lcdOutput.tft.spi.counter\[0\] vssd1 vssd1 vccd1 vccd1 net398
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8071__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4786__A_N allocation.game.controller.drawBlock.x_start\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9101__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ net152 _2642_ _2648_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__and3_1
X_5811_ _1733_ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6791_ _2601_ _2602_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5742_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__inv_2
X_8530_ _3299_ _3331_ _3865_ _3888_ _3333_ vssd1 vssd1 vccd1 vccd1 _3982_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_40_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8461_ _3297_ _3871_ vssd1 vssd1 vccd1 vccd1 _3914_ sky130_fd_sc_hd__and2_1
X_5673_ net72 _1554_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8392_ _3478_ _3849_ _3840_ vssd1 vssd1 vccd1 vccd1 _3850_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4624_ allocation.game.controller.drawBlock.x_end\[4\] allocation.game.controller.drawBlock.x_start\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7412_ net55 _3024_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__nand2_1
X_4555_ _4457_ allocation.game.controller.v\[1\] vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7343_ allocation.game.lcdOutput.tft.remainingDelayTicks\[1\] allocation.game.lcdOutput.tft.remainingDelayTicks\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4486_ allocation.game.controller.init_module.idx\[2\] vssd1 vssd1 vccd1 vccd1 _0426_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_41_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7274_ allocation.game.controller.init_module.delay_counter\[5\] _2937_ net123 vssd1
+ vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9013_ net255 vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6225_ _1052_ _2149_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__xnor2_1
X_6156_ _2019_ _2067_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__xor2_1
X_5107_ _1031_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout188_X net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6087_ _2009_ _2010_ _2011_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__and3_1
X_5038_ _0961_ _0962_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Left_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6989_ _2729_ net92 _2728_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__and3b_1
X_8728_ _2274_ _3594_ vssd1 vssd1 vccd1 vccd1 _4179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8659_ _4100_ _4101_ vssd1 vssd1 vccd1 vccd1 _4110_ sky130_fd_sc_hd__nand2_1
X_9534__315 vssd1 vssd1 vccd1 vccd1 _9534__315/HI net315 sky130_fd_sc_hd__conb_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__clkbuf_4
Xoutput8 net8 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__clkbuf_4
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9036__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6010_ _1932_ _1934_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__nand2_1
X_7961_ net137 _3473_ vssd1 vssd1 vccd1 vccd1 _3474_ sky130_fd_sc_hd__nor2_1
XANTENNA__8704__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7892_ net94 _3425_ _3426_ net108 allocation.game.controller.drawBlock.counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a32o_1
X_6912_ allocation.game.cactusDist.clock_div_inst0.counter\[5\] _2681_ vssd1 vssd1
+ vccd1 vccd1 _2683_ sky130_fd_sc_hd__and2_1
XANTENNA__8367__A1 _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6843_ allocation.game.cactus2size.clock_div_inst0.counter\[10\] _2634_ _2636_ vssd1
+ vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6774_ net160 _2591_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8513_ _3964_ vssd1 vssd1 vccd1 vccd1 _3965_ sky130_fd_sc_hd__inv_2
X_5725_ net65 _1594_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__xnor2_1
X_9493_ clknet_leaf_16_clk _0393_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.r_cactus
+ sky130_fd_sc_hd__dfxtp_1
X_5656_ _0784_ _1580_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8444_ _3334_ _3867_ _3896_ vssd1 vssd1 vccd1 vccd1 _3897_ sky130_fd_sc_hd__o21a_1
X_4607_ _0538_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoY\[4\] sky130_fd_sc_hd__inv_2
XANTENNA__7342__A2 _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8375_ _3829_ _3830_ _3836_ net197 allocation.game.controller.drawBlock.y_end\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__o32a_1
XFILLER_0_5_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5587_ _1485_ _1510_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5127__X _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4538_ allocation.game.dinoJump.count\[3\] allocation.game.dinoJump.count\[2\] allocation.game.dinoJump.count\[5\]
+ allocation.game.dinoJump.count\[4\] vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__or4_1
X_7326_ net221 allocation.game.cactusMove.drawDoneCactus net151 _2313_ vssd1 vssd1
+ vccd1 vccd1 _2972_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout103_X net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7257_ _2821_ _2926_ vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__and2_1
X_4469_ net272 vssd1 vssd1 vccd1 vccd1 _4458_ sky130_fd_sc_hd__inv_2
X_6208_ _1173_ _1227_ _2131_ _1171_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7188_ net148 _2868_ _2874_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__and3_1
XANTENNA__9059__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6139_ _2049_ _2051_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8358__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6134__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6044__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _1432_ _1433_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6490_ net92 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5441_ _1341_ _1363_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__a21oi_1
X_8160_ net473 net206 _3651_ _3657_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__o22a_1
X_5372_ _0975_ _1201_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7111_ allocation.game.controller.init_module.delay_counter\[22\] allocation.game.controller.init_module.delay_counter\[23\]
+ _2821_ _2822_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__or4_1
XANTENNA__7088__A1 allocation.game.controller.drawBlock.y_end\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8091_ _0685_ _3594_ vssd1 vssd1 vccd1 vccd1 _3595_ sky130_fd_sc_hd__nand2b_2
Xfanout107 _3479_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_2
X_7042_ allocation.game.controller.drawBlock.idx\[3\] allocation.game.controller.drawBlock.idx\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__or2_1
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout129 allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1 vccd1
+ net129 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4946__B _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8588__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8588__B2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9351__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8993_ _0655_ net52 _4440_ _4441_ vssd1 vssd1 vccd1 vccd1 _4442_ sky130_fd_sc_hd__a22o_1
X_7944_ net369 _0695_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout265_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7875_ net94 _3413_ _3414_ net108 allocation.game.controller.drawBlock.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6826_ net443 _2623_ net156 vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7563__A2 _2526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6757_ _2578_ _2579_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5708_ _1588_ _1589_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_21_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9476_ clknet_leaf_7_clk _0383_ net194 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.v\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_6688_ _2530_ _2531_ _2532_ _2533_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5639_ _1517_ _1562_ _1563_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__or3_1
X_8427_ net117 _3872_ vssd1 vssd1 vccd1 vccd1 _3880_ sky130_fd_sc_hd__nor2_1
X_8358_ net81 _2241_ _3819_ _3820_ vssd1 vssd1 vccd1 vccd1 _3821_ sky130_fd_sc_hd__o211a_1
X_7309_ net123 _2961_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__nor2_1
Xhold161 allocation.game.cactusMove.cactusMovement vssd1 vssd1 vccd1 vccd1 net484
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 allocation.game.controller.drawBlock.x_end\[8\] vssd1 vssd1 vccd1 vccd1 net473
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8276__B1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8289_ _3755_ vssd1 vssd1 vccd1 vccd1 _3756_ sky130_fd_sc_hd__inv_2
XANTENNA__7800__X _3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4872__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8751__A1 _3228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9224__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9374__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5990_ _1914_ _1913_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4941_ _0833_ _0865_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4872_ _0710_ net78 vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__nor2_4
X_7660_ allocation.game.lcdOutput.framebufferIndex\[8\] net58 vssd1 vssd1 vccd1 vccd1
+ _3222_ sky130_fd_sc_hd__xnor2_2
XANTENNA_hold86_A allocation.game.controller.drawBlock.y_start\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6611_ allocation.game.cactusMove.count\[13\] _2482_ _2484_ _2462_ vssd1 vssd1 vccd1
+ vccd1 allocation.game.cactusMove.n_count\[13\] sky130_fd_sc_hd__o211a_1
X_9330_ clknet_leaf_6_clk _0113_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7591_ _3167_ _3168_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6542_ allocation.game.dinoJump.dinoDelay\[13\] _2436_ vssd1 vssd1 vccd1 vccd1 _2437_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6473_ allocation.game.scoreCounter.clock_div.counter\[22\] allocation.game.scoreCounter.clock_div.counter\[19\]
+ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9261_ clknet_leaf_2_clk _0053_ net188 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_9192_ clknet_leaf_12_clk net354 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.tft_dc
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8212_ _0693_ _3700_ _2405_ vssd1 vssd1 vccd1 vccd1 _3701_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5424_ _1344_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__nand2_1
X_8143_ net219 _0618_ vssd1 vssd1 vccd1 vccd1 _3642_ sky130_fd_sc_hd__nand2_1
XANTENNA__7333__A _2973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5355_ _1274_ _1277_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8074_ _3565_ _3580_ _0541_ vssd1 vssd1 vccd1 vccd1 _3581_ sky130_fd_sc_hd__a21oi_1
X_5286_ _1209_ _1210_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__nand2_1
X_7025_ allocation.game.scoreCounter.bcd_tens\[6\] _2752_ allocation.game.scoreCounter.bcd_tens\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__o21ba_1
XANTENNA__4963__Y _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8976_ _3181_ _3647_ vssd1 vssd1 vccd1 vccd1 _4425_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7927_ allocation.game.controller.drawBlock.counter\[18\] _3449_ vssd1 vssd1 vccd1
+ vccd1 _3451_ sky130_fd_sc_hd__or2_1
X_7858_ allocation.game.controller.drawBlock.idx\[4\] _2762_ _2769_ _2785_ vssd1 vssd1
+ vccd1 vccd1 _3404_ sky130_fd_sc_hd__and4b_1
X_6809_ net352 _2611_ _2613_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7789_ _3319_ _3331_ _3350_ _3321_ vssd1 vssd1 vccd1 vccd1 _3351_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9247__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9528_ net322 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_19_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9459_ clknet_leaf_17_clk _0366_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__9397__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout83_X net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5710__A1 net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5140_ _0821_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5071_ _0950_ _0995_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4783__Y _0708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8830_ net268 net264 _3770_ net261 vssd1 vssd1 vccd1 vccd1 _4280_ sky130_fd_sc_hd__a31o_1
XANTENNA__5401__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5973_ _1897_ _1896_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8761_ _3874_ _4209_ _4210_ vssd1 vssd1 vccd1 vccd1 _4211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4924_ _0847_ _0848_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__and2_1
X_7712_ _3258_ _3273_ vssd1 vssd1 vccd1 vccd1 _3274_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_47_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9521__306 vssd1 vssd1 vccd1 vccd1 _9521__306/HI net306 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_23_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8692_ net76 _4123_ _4124_ _4131_ vssd1 vssd1 vccd1 vccd1 _4143_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_47_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4855_ _0774_ _0779_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7643_ allocation.game.lcdOutput.framebufferIndex\[9\] _3193_ _3203_ _3204_ vssd1
+ vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__and4_1
X_4786_ allocation.game.controller.drawBlock.x_start\[0\] allocation.game.controller.drawBlock.x_end\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__and2b_4
X_7574_ allocation.game.cactus1size.lfsr1\[0\] _3158_ net143 vssd1 vssd1 vccd1 vccd1
+ _3159_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout130_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9313_ clknet_leaf_5_clk _0105_ net173 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6525_ _2425_ _2426_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9244_ clknet_leaf_4_clk _0260_ net185 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.lfsr2\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_6456_ net225 net223 vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__and2_2
XFILLER_0_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6387_ net226 _0619_ allocation.game.cactusMove.pixel\[5\] vssd1 vssd1 vccd1 vccd1
+ _2311_ sky130_fd_sc_hd__o21a_1
X_5407_ _0751_ _0949_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9175_ clknet_leaf_16_clk _0237_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.initSeqCounter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_8126_ net112 _3614_ vssd1 vssd1 vccd1 vccd1 _3626_ sky130_fd_sc_hd__nor2_1
X_5338_ _1253_ _1256_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__a21o_1
X_8057_ _0485_ _0503_ _3519_ _0483_ vssd1 vssd1 vccd1 vccd1 _3565_ sky130_fd_sc_hd__a31o_1
XANTENNA__4974__X _0899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5269_ _1191_ _1192_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__xnor2_1
X_7008_ allocation.game.bcd_ones\[1\] _0450_ allocation.game.bcd_ones\[3\] allocation.game.bcd_ones\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8959_ _4396_ _4397_ _4407_ vssd1 vssd1 vccd1 vccd1 _4408_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_41_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6142__A _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4565__A_N allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9412__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload6_A clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _0551_ _0569_ _0550_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_42_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4571_ net262 net231 vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__xnor2_4
X_6310_ allocation.game.controller.drawBlock.state\[2\] _0606_ vssd1 vssd1 vccd1 vccd1
+ _2235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7290_ allocation.game.controller.init_module.delay_counter\[11\] allocation.game.controller.init_module.delay_counter\[10\]
+ _2946_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6241_ _1480_ _2122_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6172_ _2080_ _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5123_ _1045_ _1046_ _1047_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__nor3_1
XFILLER_0_23_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_17_clk_X clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7987__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9092__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5054_ _0798_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5131__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8813_ net38 _4250_ vssd1 vssd1 vccd1 vccd1 _4263_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8744_ _4186_ _4193_ _4184_ vssd1 vssd1 vccd1 vccd1 _4195_ sky130_fd_sc_hd__o21ba_1
X_5956_ _1861_ _1862_ _1818_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__a21oi_1
X_4907_ _0779_ _0800_ _0802_ _0777_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__o2bb2a_1
X_5887_ _1769_ _1771_ _1770_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__a21o_1
X_8675_ net89 _4125_ vssd1 vssd1 vccd1 vccd1 _4126_ sky130_fd_sc_hd__or2_1
X_4838_ _0709_ _0761_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__nand2_4
X_7626_ allocation.game.lcdOutput.framebufferIndex\[16\] allocation.game.lcdOutput.framebufferIndex\[14\]
+ allocation.game.lcdOutput.framebufferIndex\[12\] allocation.game.lcdOutput.framebufferIndex\[13\]
+ allocation.game.lcdOutput.framebufferIndex\[15\] vssd1 vssd1 vccd1 vccd1 _3188_
+ sky130_fd_sc_hd__a41o_1
X_4769_ allocation.game.controller.init_module.state\[1\] allocation.game.controller.init_module.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9046__Q allocation.game.collision.dinoY\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7557_ net340 allocation.game.lcdOutput.tft.spi.data\[4\] net256 vssd1 vssd1 vccd1
+ vccd1 _0245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6508_ allocation.game.dinoJump.dinoDelay\[0\] _2415_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[0\]
+ sky130_fd_sc_hd__and2b_1
X_7488_ _3077_ _3094_ _3083_ _3022_ vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__o2bb2a_1
X_6439_ _2361_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__inv_2
X_9227_ clknet_leaf_0_clk _0020_ net178 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9158_ clknet_leaf_18_clk _0220_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.state\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8109_ allocation.game.controller.state\[2\] _3609_ _3610_ net239 net281 vssd1 vssd1
+ vccd1 vccd1 _3611_ sky130_fd_sc_hd__a221o_1
X_9089_ clknet_leaf_14_clk _0185_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__9435__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 _0243_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 allocation.game.lcdOutput.tft.spi.data\[4\] vssd1 vssd1 vccd1 vccd1 net355
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 allocation.game.cactusDist.clock_div_inst1.counter\[13\] vssd1 vssd1 vccd1
+ vccd1 net333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold65 allocation.game.scoreCounter.clock_div.counter\[20\] vssd1 vssd1 vccd1 vccd1
+ net388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 allocation.game.cactus1size.clock_div_inst0.clk1 vssd1 vssd1 vccd1 vccd1 net377
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 allocation.game.lcdOutput.tft.remainingDelayTicks\[21\] vssd1 vssd1 vccd1
+ vccd1 net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 allocation.game.controller.init_module.delay_counter\[18\] vssd1 vssd1 vccd1
+ vccd1 net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 allocation.game.scoreCounter.bcd_tens\[4\] vssd1 vssd1 vccd1 vccd1 net421
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 allocation.game.controller.drawBlock.x_start\[6\] vssd1 vssd1 vccd1 vccd1
+ net410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8927__A1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout46_X net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5810_ _0777_ _0903_ _1733_ _1734_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__nand4_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6790_ net458 _2600_ net153 vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_44_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5741_ _1663_ _1664_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__xor2_1
X_8460_ _3889_ _3895_ _3912_ _3366_ vssd1 vssd1 vccd1 vccd1 _3913_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7411_ allocation.game.lcdOutput.tft.state\[0\] _3030_ vssd1 vssd1 vccd1 vccd1 _3032_
+ sky130_fd_sc_hd__nand2_1
X_5672_ _1596_ net82 vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__and2b_1
XANTENNA__9308__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8391_ allocation.game.controller.v\[3\] _3476_ vssd1 vssd1 vccd1 vccd1 _3849_ sky130_fd_sc_hd__and2_1
X_4623_ allocation.game.controller.drawBlock.x_start\[4\] allocation.game.controller.drawBlock.x_end\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4554_ net276 allocation.game.controller.v\[2\] vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__nand2_1
X_7342_ allocation.game.cactusHeight1\[5\] _2976_ _2978_ _2981_ vssd1 vssd1 vccd1
+ vccd1 _0201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7273_ _2937_ _2938_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__nor2_1
X_4485_ allocation.game.controller.init_module.idx\[1\] vssd1 vssd1 vccd1 vccd1 _0425_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6224_ _1008_ _2148_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9012_ net255 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6155_ _2078_ _2079_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__nand2_1
XANTENNA__8082__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5106_ _0990_ _1029_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__xor2_2
X_6086_ _1972_ _1984_ _2008_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__a21o_1
X_5037_ _0958_ _0960_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5796__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6988_ allocation.game.scoreCounter.clock_div.counter\[21\] allocation.game.scoreCounter.clock_div.counter\[20\]
+ _2725_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__and3_1
X_8727_ _4152_ _4170_ _4177_ _3996_ vssd1 vssd1 vccd1 vccd1 _4178_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5939_ _0800_ _0895_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8658_ _4107_ _4108_ vssd1 vssd1 vccd1 vccd1 _4109_ sky130_fd_sc_hd__nor2_1
X_8589_ net96 _4034_ _4037_ vssd1 vssd1 vccd1 vccd1 _4040_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7609_ net232 allocation.game.game.score\[0\] _3177_ vssd1 vssd1 vccd1 vccd1 _0273_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_47_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__clkbuf_4
Xoutput9 net9 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__clkbuf_4
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8347__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4875__A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6330__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6075__B1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7960_ _4456_ _4457_ vssd1 vssd1 vccd1 vccd1 _3473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4791__Y _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7891_ allocation.game.controller.drawBlock.counter\[7\] _3423_ vssd1 vssd1 vccd1
+ vccd1 _3426_ sky130_fd_sc_hd__or2_1
X_6911_ _2681_ _2682_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6842_ allocation.game.cactus2size.clock_div_inst0.counter\[10\] _2634_ net160 vssd1
+ vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9130__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6773_ _2590_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8512_ _3866_ _3887_ _3331_ _3373_ vssd1 vssd1 vccd1 vccd1 _3964_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5724_ _1634_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nand2_1
X_9492_ clknet_leaf_15_clk _0392_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.r_dino
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5655_ _1539_ _1541_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__xnor2_1
X_8443_ _3335_ _3868_ _3333_ vssd1 vssd1 vccd1 vccd1 _3896_ sky130_fd_sc_hd__a21o_1
XANTENNA__9280__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8374_ _3593_ _3834_ _3835_ vssd1 vssd1 vccd1 vccd1 _3836_ sky130_fd_sc_hd__or3b_1
X_4606_ net106 _0537_ _0535_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7325_ _0427_ _2970_ _2971_ net122 vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5586_ _1485_ _1510_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__nand2_1
X_4537_ allocation.game.dinoJump.count\[16\] allocation.game.dinoJump.count\[19\]
+ allocation.game.dinoJump.count\[20\] _0474_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7256_ allocation.game.controller.init_module.state\[1\] allocation.game.controller.init_module.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__and2b_1
XANTENNA__4966__Y _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4468_ net278 vssd1 vssd1 vccd1 vccd1 _4457_ sky130_fd_sc_hd__inv_2
X_6207_ _1173_ _1227_ _2131_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__nand3_1
X_7187_ allocation.game.dinoJump.count\[3\] allocation.game.dinoJump.count\[5\] allocation.game.dinoJump.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6138_ _2062_ _2061_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6069_ _1990_ _1992_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6134__B _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8597__A2 _3609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9153__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8805__A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5280__A1 _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6060__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5440_ _1315_ _1364_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5371_ _1293_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7110_ allocation.game.controller.init_module.delay_counter\[21\] allocation.game.controller.init_module.delay_counter\[20\]
+ allocation.game.controller.init_module.delay_counter\[19\] allocation.game.controller.init_module.delay_counter\[18\]
+ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8090_ net257 net164 vssd1 vssd1 vccd1 vccd1 _3594_ sky130_fd_sc_hd__nand2_1
X_7041_ allocation.game.controller.drawBlock.idx\[0\] allocation.game.controller.drawBlock.idx\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__nand2_1
Xfanout119 _3181_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_2
Xfanout108 net109 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
X_8992_ _0645_ net49 vssd1 vssd1 vccd1 vccd1 _4441_ sky130_fd_sc_hd__nand2_1
X_7943_ net384 _0695_ _2826_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4962__B _0708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8434__B net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout258_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7874_ allocation.game.controller.drawBlock.counter\[0\] allocation.game.controller.drawBlock.counter\[1\]
+ allocation.game.controller.drawBlock.counter\[2\] vssd1 vssd1 vccd1 vccd1 _3414_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout160_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6825_ allocation.game.cactus2size.clock_div_inst0.counter\[3\] allocation.game.cactus2size.clock_div_inst0.counter\[4\]
+ _2622_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_34_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6756_ net436 _2577_ net154 vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5707_ _1631_ _1630_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_21_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9475_ clknet_leaf_7_clk _0382_ net194 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.v\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6687_ allocation.game.cactus1size.clock_div_inst1.counter\[11\] allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ allocation.game.cactus1size.clock_div_inst1.counter\[13\] allocation.game.cactus1size.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5638_ _1513_ _1514_ _1516_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__a21oi_1
X_8426_ net117 net70 _3870_ vssd1 vssd1 vccd1 vccd1 _3879_ sky130_fd_sc_hd__or3_1
X_8357_ _2293_ net100 _2411_ _3562_ _3633_ vssd1 vssd1 vccd1 vccd1 _3820_ sky130_fd_sc_hd__o221a_1
XANTENNA__9026__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5569_ _0770_ _0888_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__nor2_1
Xhold151 allocation.game.controller.init_module.delay_counter\[11\] vssd1 vssd1 vccd1
+ vccd1 net474 sky130_fd_sc_hd__dlygate4sd3_1
X_7308_ allocation.game.controller.init_module.delay_counter\[17\] allocation.game.controller.init_module.delay_counter\[16\]
+ _2957_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__and3_1
XANTENNA__8276__A1 allocation.game.controller.state\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 allocation.game.dinoJump.dinoDelay\[14\] vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 allocation.game.cactusDist.clock_div_inst1.counter\[9\] vssd1 vssd1 vccd1
+ vccd1 net485 sky130_fd_sc_hd__dlygate4sd3_1
X_8288_ _0495_ _0500_ vssd1 vssd1 vccd1 vccd1 _3755_ sky130_fd_sc_hd__nor2_1
XANTENNA__8028__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7239_ net148 _0471_ _2910_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__and3_1
XANTENNA__9176__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout73_A _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4872__B net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8267__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7242__A2 _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4782__B _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4940_ _0772_ _0830_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4871_ _0768_ _0776_ _0575_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__a21o_1
X_6610_ allocation.game.cactusMove.count\[13\] _2482_ vssd1 vssd1 vccd1 vccd1 _2484_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7590_ allocation.game.cactus2size.clock_div_inst1.clk1 allocation.game.cactus2size.lfsr2\[0\]
+ allocation.game.cactus2size.lfsr2\[1\] net144 vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__a31o_1
XANTENNA__9049__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6541_ _2436_ _2415_ _2435_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[12\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_15_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6472_ allocation.game.scoreCounter.clock_div.counter\[21\] allocation.game.scoreCounter.clock_div.counter\[20\]
+ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9260_ clknet_leaf_2_clk _0048_ net181 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_8211_ net89 _0692_ vssd1 vssd1 vccd1 vccd1 _3700_ sky130_fd_sc_hd__nand2_1
X_9191_ clknet_leaf_15_clk net423 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.idle
+ sky130_fd_sc_hd__dfxtp_2
X_5423_ _0938_ _1201_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__or2_1
X_8142_ _3639_ _3640_ allocation.game.controller.state\[7\] vssd1 vssd1 vccd1 vccd1
+ _3641_ sky130_fd_sc_hd__o21a_1
X_5354_ _1225_ _1278_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8073_ _4459_ net231 vssd1 vssd1 vccd1 vccd1 _3580_ sky130_fd_sc_hd__or2_1
XANTENNA__4676__C _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5285_ net60 _1186_ _1189_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7024_ allocation.game.scoreCounter.bcd_tens\[5\] allocation.game.scoreCounter.bcd_tens\[2\]
+ allocation.game.scoreCounter.bcd_tens\[4\] vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5244__A1 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8164__B net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8975_ _0651_ net76 net69 _0660_ vssd1 vssd1 vccd1 vccd1 _4424_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_2_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout163_X net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8981__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7926_ _3449_ _3450_ allocation.game.controller.drawBlock.counter\[17\] net109 vssd1
+ vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__a2bb2o_1
X_7857_ _3402_ _3403_ _0443_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6808_ net352 _2611_ net154 vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__o21ai_1
X_7788_ _3302_ _3347_ vssd1 vssd1 vccd1 vccd1 _3350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6739_ allocation.game.cactus1size.clock_div_inst0.counter\[3\] _2566_ net154 vssd1
+ vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9527_ net321 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
X_9458_ clknet_leaf_18_clk _0365_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_8409_ net43 _3276_ _3356_ net34 vssd1 vssd1 vccd1 vccd1 _3862_ sky130_fd_sc_hd__o31a_1
X_9389_ clknet_leaf_13_clk _0299_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.idx\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout76_X net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__B _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8090__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7932__B1 _3410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout90 _2414_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
XFILLER_0_49_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9341__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9491__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5070_ _0993_ _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__nor2_1
X_5972_ _1843_ _1848_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__xnor2_1
X_8760_ net48 _3308_ _3930_ vssd1 vssd1 vccd1 vccd1 _4210_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4923_ _0788_ _0841_ _0846_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__or3_1
X_7711_ _3252_ _3257_ vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8691_ _3237_ _3595_ _4093_ _4141_ _4140_ vssd1 vssd1 vccd1 vccd1 _4142_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_47_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4854_ _0710_ _0778_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__nor2_2
X_7642_ allocation.game.lcdOutput.framebufferIndex\[10\] _3198_ _3201_ vssd1 vssd1
+ vccd1 vccd1 _3204_ sky130_fd_sc_hd__o21ba_1
XANTENNA__7923__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4785_ _0707_ _0708_ _0605_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__a21o_4
XANTENNA__7328__B net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7573_ net377 allocation.game.cactus1size.lfsr1\[1\] vssd1 vssd1 vccd1 vccd1 _3158_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6524_ allocation.game.dinoJump.dinoDelay\[6\] _2423_ _2415_ vssd1 vssd1 vccd1 vccd1
+ _2426_ sky130_fd_sc_hd__o21ai_1
X_9312_ clknet_leaf_2_clk _0272_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.clk1
+ sky130_fd_sc_hd__dfxtp_1
X_9243_ clknet_leaf_3_clk _0259_ net193 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.lfsr2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6455_ _2373_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4968__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5406_ _0939_ _1179_ _0940_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__a21o_1
X_6386_ _2267_ _2296_ _2309_ _2304_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__a31o_1
X_9174_ clknet_leaf_19_clk _0236_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.initSeqCounter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_8125_ net408 net207 _3625_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__o21a_1
X_5337_ _1260_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8056_ net267 _3520_ _3562_ vssd1 vssd1 vccd1 vccd1 _3564_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5268_ _1174_ _1190_ _1192_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__and3_1
X_7007_ _0450_ allocation.game.bcd_ones\[2\] _2739_ _2742_ vssd1 vssd1 vccd1 vccd1
+ net13 sky130_fd_sc_hd__a31oi_1
X_5199_ _1121_ _1123_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__and2b_1
X_8958_ _4399_ _4406_ _4400_ vssd1 vssd1 vccd1 vccd1 _4407_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9214__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7909_ net95 _3437_ _3438_ net109 allocation.game.controller.drawBlock.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8889_ net259 _3261_ _3264_ net261 _4338_ vssd1 vssd1 vccd1 vccd1 _4339_ sky130_fd_sc_hd__o221ai_1
XANTENNA__9364__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6142__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4878__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8890__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout280 allocation.game.collision.dinoY\[0\] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4570_ net267 allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_42_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8881__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6240_ _1424_ _2123_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__nor2_1
X_6171_ _2087_ _2095_ _2088_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__o21a_1
XANTENNA__9088__RESET_B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5122_ _1009_ _1043_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__and2_1
XANTENNA__9237__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5053_ _0806_ _0846_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8812_ net44 _4261_ vssd1 vssd1 vccd1 vccd1 _4262_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9387__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5955_ _1864_ _1877_ _1878_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__nand3_1
X_8743_ _4184_ _4186_ _4192_ vssd1 vssd1 vccd1 vccd1 _4194_ sky130_fd_sc_hd__or3_1
X_4906_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8674_ _0673_ _4122_ vssd1 vssd1 vccd1 vccd1 _4125_ sky130_fd_sc_hd__nor2_1
X_5886_ _1798_ _1799_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__xnor2_1
X_4837_ _0737_ _0755_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7625_ _3179_ _3183_ vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__nor2_1
X_4768_ allocation.game.controller.block_done allocation.game.controller.state\[7\]
+ _0684_ _0694_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a211o_1
X_7556_ net335 allocation.game.lcdOutput.tft.spi.data\[3\] net256 vssd1 vssd1 vccd1
+ vccd1 _0244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4699_ _0618_ _0624_ allocation.game.controller.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _0627_ sky130_fd_sc_hd__o21ai_2
X_6507_ _0461_ _2414_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__and2b_2
X_7487_ _3045_ _3046_ _3094_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__or3_1
X_6438_ _2334_ _2349_ _2338_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__o21a_1
XANTENNA__8872__A1 _0401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9226_ clknet_leaf_2_clk _0256_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.clk1
+ sky130_fd_sc_hd__dfxtp_1
X_9157_ clknet_leaf_12_clk _0219_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.color\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8108_ _0612_ _2518_ vssd1 vssd1 vccd1 vccd1 _3610_ sky130_fd_sc_hd__nand2_1
X_6369_ allocation.game.cactusHeight1\[5\] _2291_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__or2_1
X_9088_ clknet_leaf_14_clk _0184_ net215 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold22 allocation.game.lcdOutput.tft.spi.data\[5\] vssd1 vssd1 vccd1 vccd1 net345
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 allocation.game.cactus1size.clock_div_inst0.counter\[13\] vssd1 vssd1 vccd1
+ vccd1 net334 sky130_fd_sc_hd__dlygate4sd3_1
X_8039_ _3531_ _3546_ vssd1 vssd1 vccd1 vccd1 _3548_ sky130_fd_sc_hd__nand2_1
Xhold55 allocation.game.scoreCounter.clock_div.counter\[23\] vssd1 vssd1 vccd1 vccd1
+ net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 allocation.game.lcdOutput.tft.spi.data\[3\] vssd1 vssd1 vccd1 vccd1 net356
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 allocation.game.lcdOutput.tft.spi.data\[7\] vssd1 vssd1 vccd1 vccd1 net367
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 allocation.game.controller.drawBlock.y_start\[2\] vssd1 vssd1 vccd1 vccd1
+ net400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 allocation.game.controller.drawBlock.x_end\[2\] vssd1 vssd1 vccd1 vccd1 net389
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 allocation.game.controller.drawBlock.x_end\[6\] vssd1 vssd1 vccd1 vccd1 net411
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 allocation.game.lcdOutput.tft.spi.idle vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_27_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8615__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6626__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5740_ _1664_ _1663_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _0727_ net88 _1123_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__a21oi_1
X_7410_ allocation.game.lcdOutput.tft.state\[2\] allocation.game.lcdOutput.tft.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__or2_1
X_8390_ allocation.game.controller.v\[3\] net85 vssd1 vssd1 vccd1 vccd1 _3848_ sky130_fd_sc_hd__and2b_1
X_4622_ _0550_ _0551_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_26_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4553_ _0487_ _0489_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7341_ net486 _2975_ _2980_ _2982_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4484_ allocation.game.controller.init_module.idx\[0\] vssd1 vssd1 vccd1 vccd1 _0424_
+ sky130_fd_sc_hd__inv_2
X_7272_ net425 _2935_ net122 vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6223_ _1016_ _1021_ _1019_ _0841_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9011_ net255 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6154_ _2076_ _2077_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__nand2b_1
XANTENNA__8082__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5105_ net82 _0820_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__and3_1
X_6085_ _1874_ _1918_ _1919_ _1923_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__a31o_1
X_5036_ _0958_ _0960_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6987_ allocation.game.scoreCounter.clock_div.counter\[20\] allocation.game.scoreCounter.clock_div.counter\[19\]
+ _2724_ allocation.game.scoreCounter.clock_div.counter\[21\] vssd1 vssd1 vccd1 vccd1
+ _2728_ sky130_fd_sc_hd__a31o_1
XANTENNA__5796__B _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8726_ _4172_ _4175_ _4176_ _0669_ vssd1 vssd1 vccd1 vccd1 _4177_ sky130_fd_sc_hd__o31a_1
X_5938_ _1819_ _1861_ _1862_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5869_ _1766_ _1777_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__xor2_1
X_8657_ _4101_ _4103_ vssd1 vssd1 vccd1 vccd1 _4108_ sky130_fd_sc_hd__nand2_1
X_8588_ net67 _3621_ _4038_ net74 vssd1 vssd1 vccd1 vccd1 _4039_ sky130_fd_sc_hd__a22o_1
X_7608_ allocation.game.game.score\[0\] _2328_ _3176_ _2319_ net145 vssd1 vssd1 vccd1
+ vccd1 _3177_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9402__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7539_ allocation.game.lcdOutput.tft.state\[0\] _3031_ _3037_ _3020_ vssd1 vssd1
+ vccd1 vccd1 _3147_ sky130_fd_sc_hd__o211a_1
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
X_9209_ _0147_ _0406_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6608__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6148__A _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_16_clk_X clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9082__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6311__A2 allocation.game.controller.drawBlock.state\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6075__B2 _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6075__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5897__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7890_ allocation.game.controller.drawBlock.counter\[7\] _3423_ vssd1 vssd1 vccd1
+ vccd1 _3425_ sky130_fd_sc_hd__nand2_1
X_6910_ allocation.game.cactusDist.clock_div_inst0.counter\[4\] _2679_ net155 vssd1
+ vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6841_ _2634_ _2635_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8511_ _3330_ _3962_ vssd1 vssd1 vccd1 vccd1 _3963_ sky130_fd_sc_hd__nand2_1
X_6772_ _2587_ _2588_ _2589_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__or3_1
XANTENNA__9425__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5723_ _1634_ _1646_ _1647_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__nand3_1
X_9491_ clknet_leaf_20_clk _0391_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.r_cloud
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5654_ _1542_ _1543_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__xor2_1
X_8442_ _3289_ _3291_ _3304_ _3868_ vssd1 vssd1 vccd1 vccd1 _3895_ sky130_fd_sc_hd__a22oi_2
X_4605_ _0505_ _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__nor2_1
X_8373_ _2292_ net100 _2411_ _3578_ _3633_ vssd1 vssd1 vccd1 vccd1 _3835_ sky130_fd_sc_hd__o221a_1
X_7324_ _0427_ _2970_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__nand2_1
XANTENNA__4679__C net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5585_ net65 _1458_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__xor2_1
X_4536_ allocation.game.dinoJump.count\[13\] allocation.game.dinoJump.count\[15\]
+ allocation.game.dinoJump.count\[14\] allocation.game.dinoJump.count\[12\] vssd1
+ vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__or4b_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7255_ _4459_ allocation.game.dinoJump.next_dinoY\[6\] _2915_ _2925_ vssd1 vssd1
+ vccd1 vccd1 _0171_ sky130_fd_sc_hd__a211o_1
X_4467_ net280 vssd1 vssd1 vccd1 vccd1 _4456_ sky130_fd_sc_hd__inv_2
XANTENNA__4976__A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7186_ allocation.game.dinoJump.count\[4\] _2870_ allocation.game.dinoJump.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__a21oi_1
X_6206_ _1282_ _1327_ _2129_ _1280_ _1230_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__a311o_1
X_6137_ _1858_ _2029_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__xnor2_1
X_6068_ net103 net124 vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__nor2_1
X_5019_ _0752_ _0942_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8709_ net120 _4154_ vssd1 vssd1 vccd1 vccd1 _4160_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5370_ _1242_ _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4796__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7040_ _0443_ _0444_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout109 _3409_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8991_ net257 _3249_ _4168_ vssd1 vssd1 vccd1 vccd1 _4440_ sky130_fd_sc_hd__a21bo_1
X_7942_ allocation.game.controller.init_module.idx\[0\] allocation.game.controller.init_module.idx\[1\]
+ _2825_ _0398_ allocation.game.controller.init_module.idx\[2\] vssd1 vssd1 vccd1
+ vccd1 _0324_ sky130_fd_sc_hd__a311o_1
XFILLER_0_37_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5420__A _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7873_ allocation.game.controller.drawBlock.counter\[0\] allocation.game.controller.drawBlock.counter\[1\]
+ allocation.game.controller.drawBlock.counter\[2\] vssd1 vssd1 vccd1 vccd1 _3413_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout153_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6824_ _2623_ _2624_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6755_ allocation.game.cactus1size.clock_div_inst0.counter\[9\] _2577_ vssd1 vssd1
+ vccd1 vccd1 _2578_ sky130_fd_sc_hd__and2_1
X_9474_ clknet_leaf_7_clk _0381_ net194 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.v\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_5706_ _1027_ _1618_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6686_ allocation.game.cactus1size.clock_div_inst1.counter\[7\] allocation.game.cactus1size.clock_div_inst1.counter\[6\]
+ allocation.game.cactus1size.clock_div_inst1.counter\[9\] allocation.game.cactus1size.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__or4_1
X_8425_ net127 net45 _3279_ _3271_ vssd1 vssd1 vccd1 vccd1 _3878_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_21_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5637_ _1533_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__nand2_1
X_8356_ _3479_ _3818_ net244 vssd1 vssd1 vccd1 vccd1 _3819_ sky130_fd_sc_hd__o21ai_1
X_5568_ _0918_ _1447_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__xor2_1
X_7307_ net460 _2957_ _2960_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8287_ net277 net135 _3514_ _3753_ vssd1 vssd1 vccd1 vccd1 _3754_ sky130_fd_sc_hd__o211a_1
Xhold130 allocation.game.cactus1size.clock_div_inst1.counter\[12\] vssd1 vssd1 vccd1
+ vccd1 net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 allocation.game.dinoJump.dinoDelay\[10\] vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ allocation.game.dinoJump.dinoDelay\[7\] allocation.game.dinoJump.dinoDelay\[6\]
+ allocation.game.dinoJump.dinoDelay\[9\] allocation.game.dinoJump.dinoDelay\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__nand4_1
Xhold141 allocation.game.cactusDist.clock_div_inst1.counter\[3\] vssd1 vssd1 vccd1
+ vccd1 net464 sky130_fd_sc_hd__dlygate4sd3_1
X_7238_ _2910_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__inv_2
Xhold163 allocation.game.cactusHeight1\[4\] vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _1422_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__nor2_1
X_7169_ allocation.game.lcdOutput.tft.spi.internalSck net4 allocation.game.lcdOutput.tft.spi.cs
+ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__and3_1
XANTENNA__8028__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout66_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6211__A1 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9120__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7720__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9512__297 vssd1 vssd1 vccd1 vccd1 _9512__297/HI net297 sky130_fd_sc_hd__conb_1
XANTENNA__8975__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9270__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6450__B2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8727__B1 _3996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4870_ _0793_ _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6540_ allocation.game.dinoJump.dinoDelay\[11\] allocation.game.dinoJump.dinoDelay\[12\]
+ _2432_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
X_6471_ net146 _2359_ _2384_ _2369_ allocation.game.scoreCounter.bcd_tens\[3\] vssd1
+ vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a32o_1
XANTENNA__4797__Y _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8210_ _0680_ _3647_ _3698_ vssd1 vssd1 vccd1 vccd1 _3699_ sky130_fd_sc_hd__o21a_1
X_9190_ clknet_leaf_15_clk _0252_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_5422_ _1197_ _1346_ _1345_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8141_ _0673_ _0690_ vssd1 vssd1 vccd1 vccd1 _3640_ sky130_fd_sc_hd__nor2_1
X_5353_ net62 _1224_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8072_ _3564_ _3578_ vssd1 vssd1 vccd1 vccd1 _3579_ sky130_fd_sc_hd__xor2_1
X_5284_ _1186_ _1189_ net60 vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7023_ _0439_ allocation.game.scoreCounter.bcd_tens\[4\] _2751_ allocation.game.scoreCounter.bcd_tens\[2\]
+ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__a211o_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8974_ _2241_ net37 _3276_ _2242_ _4422_ vssd1 vssd1 vccd1 vccd1 _4423_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout270_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7925_ allocation.game.controller.drawBlock.counter\[17\] _3447_ net95 vssd1 vssd1
+ vccd1 vccd1 _3450_ sky130_fd_sc_hd__o21ai_1
X_7856_ allocation.game.controller.drawBlock.state\[3\] _3402_ vssd1 vssd1 vccd1 vccd1
+ _3403_ sky130_fd_sc_hd__nor2_1
X_6807_ _2611_ _2612_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4999_ net64 _0923_ _0893_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__a21oi_4
X_9526_ net311 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
X_7787_ _3323_ _3348_ _3346_ vssd1 vssd1 vccd1 vccd1 _3349_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6738_ allocation.game.cactus1size.clock_div_inst0.counter\[3\] _2566_ vssd1 vssd1
+ vccd1 vccd1 _2567_ sky130_fd_sc_hd__and2_1
X_6669_ net151 _2461_ _2519_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__and3_1
X_9457_ clknet_leaf_18_clk _0364_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9388_ clknet_leaf_14_clk _0298_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.idx\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8408_ _3311_ _3362_ _3359_ _3271_ vssd1 vssd1 vccd1 vccd1 _3861_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8339_ net107 _3802_ net244 vssd1 vssd1 vccd1 vccd1 _3803_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9293__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout69_X net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4994__A1 _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8185__B2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout91 net93 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
Xfanout80 _0717_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7715__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5889__B net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
X_5971_ _1893_ _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__nand2_1
X_4922_ _0841_ _0846_ _0788_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7449__X _3066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7710_ net39 net35 vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__nand2_1
X_8690_ net164 net49 vssd1 vssd1 vccd1 vccd1 _4141_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7641_ _3183_ _3202_ vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_47_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4853_ _0768_ _0776_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__xnor2_4
XANTENNA__7923__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4784_ _0707_ _0708_ _0605_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_7_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7572_ net377 _2562_ _3014_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9311_ clknet_leaf_2_clk _0271_ net181 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.lfsr2\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_6523_ allocation.game.dinoJump.dinoDelay\[6\] _2423_ vssd1 vssd1 vccd1 vccd1 _2425_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6454_ net230 net227 net226 vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__o21a_1
X_9242_ clknet_leaf_4_clk _0258_ net185 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.lfsr1\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5405_ _1329_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__inv_2
X_6385_ _2303_ _2308_ _2307_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9173_ clknet_leaf_19_clk _0235_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.initSeqCounter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_8124_ net243 _3614_ _3615_ _3624_ vssd1 vssd1 vccd1 vccd1 _3625_ sky130_fd_sc_hd__a31o_1
X_5336_ _1258_ _1259_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5267_ _1131_ _1147_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__xnor2_2
X_8055_ net265 _3520_ _3562_ vssd1 vssd1 vccd1 vccd1 _3563_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4984__A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7006_ _2739_ _2741_ _0450_ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__a21oi_1
X_5198_ _1064_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8957_ net68 _3673_ _4080_ _4405_ _4078_ vssd1 vssd1 vccd1 vccd1 _4406_ sky130_fd_sc_hd__o221a_1
X_7908_ allocation.game.controller.drawBlock.counter\[12\] _3434_ vssd1 vssd1 vccd1
+ vccd1 _3438_ sky130_fd_sc_hd__or2_1
X_8888_ net262 _3264_ _4307_ _4337_ vssd1 vssd1 vccd1 vccd1 _4338_ sky130_fd_sc_hd__a211o_1
X_7839_ allocation.game.cactus2size.lfsr1\[0\] allocation.game.cactus2size.lfsr2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3394_ sky130_fd_sc_hd__xor2_2
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload0 clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9496__318 vssd1 vssd1 vccd1 vccd1 net318 _9496__318/LO sky130_fd_sc_hd__conb_1
X_9509_ net294 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4878__B _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9039__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_4
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6170_ _2092_ _2094_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5121_ _1007_ _1009_ _1005_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7180__A _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5052_ _0805_ _0846_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8811_ _4242_ _4260_ vssd1 vssd1 vccd1 vccd1 _4261_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8742_ _4191_ _4192_ vssd1 vssd1 vccd1 vccd1 _4193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5954_ _1877_ _1878_ _1864_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__a21o_1
X_4905_ _0709_ net88 _0808_ _0807_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__a31oi_4
X_5885_ _1807_ _1809_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__and2b_1
X_8673_ net67 _3617_ _4123_ net76 vssd1 vssd1 vccd1 vccd1 _4124_ sky130_fd_sc_hd__a22o_1
X_4836_ _0737_ _0755_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__xor2_4
XFILLER_0_29_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7624_ allocation.game.lcdOutput.framebufferIndex\[12\] net120 _3179_ vssd1 vssd1
+ vccd1 vccd1 _3186_ sky130_fd_sc_hd__a21boi_1
X_7555_ allocation.game.lcdOutput.tft.spi.dataShift\[5\] net343 net256 vssd1 vssd1
+ vccd1 vccd1 _0243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4767_ _0690_ _0693_ allocation.game.controller.state\[7\] vssd1 vssd1 vccd1 vccd1
+ _0694_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_16_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6506_ _0464_ net106 vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__and2_1
X_4698_ _0618_ _0624_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__nor2_1
XANTENNA__4591__C1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7486_ net343 net53 _3072_ _3100_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout119_X net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6437_ _2359_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__inv_2
X_9225_ clknet_leaf_22_clk _0038_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_9156_ clknet_leaf_12_clk _0218_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.color\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_6368_ allocation.game.cactusHeight1\[5\] _2291_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__nor2_1
X_5319_ _1191_ _1243_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__nand2_1
X_8107_ _3608_ vssd1 vssd1 vccd1 vccd1 _3609_ sky130_fd_sc_hd__inv_2
XANTENNA__4894__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9087_ clknet_leaf_14_clk _0183_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold12 allocation.game.lcdOutput.tft.spi.dataShift\[4\] vssd1 vssd1 vccd1 vccd1 net335
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 allocation.game.lcdOutput.tft.spi.dataShift\[2\] vssd1 vssd1 vccd1 vccd1 net346
+ sky130_fd_sc_hd__dlygate4sd3_1
X_6299_ allocation.game.controller.drawBlock.counter\[16\] _2175_ _2178_ _2179_ _2223_
+ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__a2111o_1
XANTENNA__5603__A _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8038_ _3531_ _3546_ vssd1 vssd1 vccd1 vccd1 _3547_ sky130_fd_sc_hd__or2_1
Xhold56 allocation.game.controller.drawBlock.x_end\[7\] vssd1 vssd1 vccd1 vccd1 net379
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 allocation.game.lcdOutput.tft.spi.data\[8\] vssd1 vssd1 vccd1 vccd1 net357
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 allocation.game.lcdOutput.tft.spi.data\[0\] vssd1 vssd1 vccd1 vccd1 net368
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9480__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 allocation.game.scoreCounter.clock_div.counter\[17\] vssd1 vssd1 vccd1 vccd1
+ net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 allocation.game.controller.drawBlock.state\[1\] vssd1 vssd1 vccd1 vccd1 net412
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 allocation.game.lcdOutput.tft.state\[2\] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9331__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8633__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9481__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8312__B2 allocation.game.controller.drawBlock.y_end\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9150__RESET_B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8543__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5670_ net65 _1594_ _1593_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4621_ allocation.game.controller.drawBlock.x_end\[5\] allocation.game.controller.drawBlock.x_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__nand2b_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552_ _0487_ _0489_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__and2_1
X_7340_ allocation.game.cactusHeight1\[3\] _2976_ _2979_ _2981_ vssd1 vssd1 vccd1
+ vccd1 _0199_ sky130_fd_sc_hd__a211o_1
X_7271_ allocation.game.controller.init_module.delay_counter\[4\] allocation.game.controller.init_module.delay_counter\[3\]
+ _2933_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__and3_1
X_4483_ allocation.game.dinoJump.drawDoneDino vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6222_ _2145_ _2146_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9010_ net255 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__inv_2
XANTENNA__8067__B1 _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6153_ _2075_ _2077_ _2074_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__or3b_1
XANTENNA__5423__A _0938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9354__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5104_ _1027_ _1028_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__and2_1
X_6084_ _1972_ _1984_ _2008_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__nand3_1
X_5035_ _0864_ _0869_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8734__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6986_ net388 _2725_ _2727_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5937_ _1772_ _1812_ _1817_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__a21o_1
XANTENNA__8790__A1 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8725_ _4156_ _4161_ _4160_ _4159_ vssd1 vssd1 vccd1 vccd1 _4176_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8656_ net104 _3190_ _4106_ vssd1 vssd1 vccd1 vccd1 _4107_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5868_ _0896_ _1790_ _1791_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__nand3_1
X_7607_ allocation.game.game.score\[0\] _2320_ vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__xor2_1
X_4819_ _0724_ _0741_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__nor2_1
X_8587_ net223 _3619_ vssd1 vssd1 vccd1 vccd1 _4038_ sky130_fd_sc_hd__xnor2_1
X_5799_ _1670_ _1721_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7538_ net357 _3146_ _0233_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7469_ allocation.game.lcdOutput.tft.initSeqCounter\[0\] net249 vssd1 vssd1 vccd1
+ vccd1 _3085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_32_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
X_9208_ _0146_ _0405_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__7813__A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8628__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout96_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9139_ clknet_leaf_18_clk _0203_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6148__B _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5052__B _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout51_X net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7336__A2 _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9227__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9377__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6075__A2 _0886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8554__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6840_ net476 _2633_ net157 vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6771_ allocation.game.cactus2size.clock_div_inst1.counter\[11\] allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ allocation.game.cactus2size.clock_div_inst1.counter\[13\] allocation.game.cactus2size.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8510_ net68 _3325_ _3961_ vssd1 vssd1 vccd1 vccd1 _3962_ sky130_fd_sc_hd__or3b_1
X_5722_ _1619_ _1632_ _1633_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9490_ clknet_leaf_20_clk _0390_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.r_over
+ sky130_fd_sc_hd__dfxtp_1
X_8441_ _3321_ net70 _3893_ net118 vssd1 vssd1 vccd1 vccd1 _3894_ sky130_fd_sc_hd__o31a_1
X_5653_ _1558_ _1577_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4604_ _0487_ _0502_ _0504_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__and3_1
X_8372_ _3831_ _3832_ _3833_ _3514_ vssd1 vssd1 vccd1 vccd1 _3834_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5584_ net65 _1508_ _1506_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__a21oi_1
X_7323_ net122 _2969_ _2970_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__and3_1
X_4535_ allocation.game.dinoJump.count\[1\] allocation.game.dinoJump.count\[0\] allocation.game.dinoJump.count\[17\]
+ allocation.game.dinoJump.count\[18\] vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_15_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7254_ net261 _0513_ _2916_ _2917_ _2924_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__a221o_1
XANTENNA__4976__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4466_ net232 vssd1 vssd1 vccd1 vccd1 _4455_ sky130_fd_sc_hd__inv_2
X_7185_ net416 _2870_ _2872_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__a21oi_1
X_6205_ _1282_ _1327_ _2129_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6136_ _2059_ _2060_ _2058_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6067_ _1951_ _1991_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__nand2_1
X_5018_ _0752_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6969_ allocation.game.scoreCounter.clock_div.counter\[14\] _2715_ vssd1 vssd1 vccd1
+ vccd1 _2717_ sky130_fd_sc_hd__and2_1
XANTENNA__7808__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8708_ _3199_ _4158_ _4156_ _4150_ vssd1 vssd1 vccd1 vccd1 _4159_ sky130_fd_sc_hd__a211o_1
XANTENNA__8515__A1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8639_ _4072_ _4082_ _4089_ _4081_ vssd1 vssd1 vccd1 vccd1 _4090_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout99_X net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7254__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8093__B net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8506__A1 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9517__302 vssd1 vssd1 vccd1 vccd1 _9517__302/HI net302 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_10_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7453__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8284__A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8990_ _4430_ _4433_ _4438_ _4436_ vssd1 vssd1 vccd1 vccd1 _4439_ sky130_fd_sc_hd__a31o_1
X_7941_ allocation.game.controller.init_module.idx\[1\] _3458_ _3459_ vssd1 vssd1
+ vccd1 vccd1 _0323_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7872_ allocation.game.controller.drawBlock.counter\[0\] allocation.game.controller.drawBlock.counter\[1\]
+ _3412_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6823_ allocation.game.cactus2size.clock_div_inst0.counter\[3\] _2622_ net155 vssd1
+ vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout146_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6754_ net160 _2576_ _2577_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__nor3_1
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9473_ clknet_leaf_8_clk _0380_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_end\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_5705_ _1621_ _1629_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__nand2_1
X_6685_ allocation.game.cactus1size.clock_div_inst1.counter\[3\] allocation.game.cactus1size.clock_div_inst1.counter\[5\]
+ allocation.game.cactus1size.clock_div_inst1.counter\[4\] allocation.game.cactus1size.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__or4b_1
XFILLER_0_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5636_ _1552_ _1559_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__xnor2_1
X_8424_ net70 _3862_ _3870_ _3876_ vssd1 vssd1 vccd1 vccd1 _3877_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_21_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8355_ net139 _3560_ _3561_ _3817_ vssd1 vssd1 vccd1 vccd1 _3818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5567_ _0773_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7306_ net123 _2959_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__nor2_1
Xhold142 allocation.game.controller.init_module.delay_counter\[0\] vssd1 vssd1 vccd1
+ vccd1 net465 sky130_fd_sc_hd__dlygate4sd3_1
X_8286_ net135 _3496_ vssd1 vssd1 vccd1 vccd1 _3753_ sky130_fd_sc_hd__nand2_1
X_4518_ allocation.game.dinoJump.dinoDelay\[11\] allocation.game.dinoJump.dinoDelay\[10\]
+ allocation.game.dinoJump.dinoDelay\[13\] allocation.game.dinoJump.dinoDelay\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__or4b_1
Xhold131 allocation.game.lcdOutput.tft.remainingDelayTicks\[5\] vssd1 vssd1 vccd1
+ vccd1 net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 allocation.game.cactus2size.clock_div_inst0.counter\[4\] vssd1 vssd1 vccd1
+ vccd1 net443 sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ _1417_ _1420_ _1421_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__and3_1
Xhold153 allocation.game.cactus2size.clock_div_inst0.counter\[9\] vssd1 vssd1 vccd1
+ vccd1 net476 sky130_fd_sc_hd__dlygate4sd3_1
X_7237_ allocation.game.dinoJump.count\[19\] _2909_ vssd1 vssd1 vccd1 vccd1 _2910_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7168_ allocation.game.lcdOutput.tft.spi.cs net4 vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__and2b_1
X_7099_ allocation.game.controller.drawBlock.y_end\[6\] _2779_ _0417_ vssd1 vssd1
+ vccd1 vccd1 _2813_ sky130_fd_sc_hd__a21o_1
X_6119_ _2002_ _2004_ _2032_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__and3_1
XANTENNA__9072__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8922__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9415__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5521__A _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__A1 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8551__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9436__Q allocation.game.controller.drawBlock.x_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6470_ net146 _2385_ _2386_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a21o_1
X_5421_ _0834_ _1198_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__xnor2_1
X_8140_ _0673_ _0690_ vssd1 vssd1 vccd1 vccd1 _3639_ sky130_fd_sc_hd__and2_1
XANTENNA__7183__A _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5352_ net62 _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8071_ net259 _3560_ vssd1 vssd1 vccd1 vccd1 _3578_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7022_ allocation.game.scoreCounter.bcd_tens\[6\] allocation.game.scoreCounter.bcd_tens\[1\]
+ allocation.game.scoreCounter.bcd_tens\[0\] allocation.game.scoreCounter.bcd_tens\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__or4_1
X_5283_ _0893_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__nor2_1
XANTENNA__9095__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7630__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8966__A1 _0401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8973_ _2242_ net37 _4421_ _4420_ vssd1 vssd1 vccd1 vccd1 _4422_ sky130_fd_sc_hd__o31a_1
X_7924_ allocation.game.controller.drawBlock.counter\[17\] _3447_ vssd1 vssd1 vccd1
+ vccd1 _3449_ sky130_fd_sc_hd__and2_1
X_7855_ allocation.game.controller.drawBlock.state\[2\] allocation.game.controller.drawBlock.state\[3\]
+ _3400_ _3401_ net236 vssd1 vssd1 vccd1 vccd1 _3402_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_37_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6806_ net445 _2610_ net154 vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4998_ _0922_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__inv_2
X_9525_ net310 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_7786_ _3317_ net114 _3288_ _3347_ vssd1 vssd1 vccd1 vccd1 _3348_ sky130_fd_sc_hd__and4b_1
X_6737_ net160 _2565_ _2566_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6668_ _2520_ net407 _2515_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_pixel\[4\]
+ sky130_fd_sc_hd__mux2_1
X_9456_ clknet_leaf_18_clk _0363_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_8407_ _3842_ _3860_ _3859_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__o21ai_1
X_9387_ clknet_leaf_14_clk _0297_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.idx\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_6599_ allocation.game.cactusMove.count\[9\] _2475_ vssd1 vssd1 vccd1 vccd1 _2477_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5619_ _1543_ _1542_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8338_ net139 _3542_ _3800_ _3801_ vssd1 vssd1 vccd1 vccd1 _3802_ sky130_fd_sc_hd__a22o_1
XANTENNA__9438__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8917__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8269_ net235 _3739_ _3738_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__mux2_1
XANTENNA__8957__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4994__A2 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout92 _2404_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout81 _0683_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout70 _3370_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9104__RESET_B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7731__A _3248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7450__B _3066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5970_ _1886_ _1893_ _1894_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4921_ net88 _0771_ _0775_ _0779_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__a22o_2
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4852_ _0768_ _0776_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__xor2_4
X_7640_ allocation.game.lcdOutput.framebufferIndex\[10\] _3193_ net74 _3192_ vssd1
+ vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_47_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7571_ _0431_ net361 _2526_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__a21o_1
X_4783_ _0602_ _0604_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4907__A2_N _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9310_ clknet_leaf_3_clk _0270_ net191 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.lfsr2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_6522_ _2423_ _2424_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6453_ allocation.game.scoreCounter.bcd_tens\[1\] _2369_ _2372_ net146 vssd1 vssd1
+ vccd1 vccd1 _0013_ sky130_fd_sc_hd__a22o_1
X_9241_ clknet_leaf_3_clk _0257_ net193 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.lfsr1\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4968__C net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5404_ _1323_ _1325_ _1326_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__a21o_1
X_9172_ clknet_leaf_19_clk _0234_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.frameBufferLowNibble
+ sky130_fd_sc_hd__dfxtp_1
X_8123_ allocation.game.controller.state\[7\] _3617_ _3621_ allocation.game.controller.state\[2\]
+ _3623_ vssd1 vssd1 vccd1 vccd1 _3624_ sky130_fd_sc_hd__a221o_1
X_6384_ _2285_ _2288_ _2290_ _2306_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout109_A _3409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5335_ _1259_ _1258_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__nand2b_1
XANTENNA__8636__B1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8054_ _3560_ _3561_ vssd1 vssd1 vccd1 vccd1 _3562_ sky130_fd_sc_hd__nand2_2
XANTENNA__4984__B _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5266_ _1174_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__nand2_1
XANTENNA__6111__A1 _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7005_ allocation.game.bcd_ones\[1\] allocation.game.bcd_ones\[3\] vssd1 vssd1 vccd1
+ vccd1 _2741_ sky130_fd_sc_hd__nand2_1
X_5197_ _0809_ _0822_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__nor2_1
XANTENNA__8939__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8956_ _4017_ _4018_ _4055_ _0619_ vssd1 vssd1 vccd1 vccd1 _4405_ sky130_fd_sc_hd__a211oi_1
X_7907_ allocation.game.controller.drawBlock.counter\[12\] _3434_ vssd1 vssd1 vccd1
+ vccd1 _3437_ sky130_fd_sc_hd__nand2_1
X_8887_ _4309_ _4325_ _4306_ _4308_ vssd1 vssd1 vccd1 vccd1 _4337_ sky130_fd_sc_hd__a211oi_1
XANTENNA__9110__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7838_ allocation.game.cactus2size.lfsr1\[1\] allocation.game.cactus2size.lfsr2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3393_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7769_ net117 net96 vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__nor2_2
X_9508_ net293 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xclkload1 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9439_ clknet_leaf_11_clk _0348_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9260__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout81_X net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout282 _0608_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
Xfanout260 allocation.game.collision.dinoY\[7\] vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xfanout271 allocation.game.collision.dinoY\[4\] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7726__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8557__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5120_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__inv_2
X_5051_ net80 _0782_ _0948_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8810_ net272 _3760_ net268 vssd1 vssd1 vccd1 vccd1 _4260_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9133__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8741_ net96 _4185_ _4190_ _3200_ vssd1 vssd1 vccd1 vccd1 _4192_ sky130_fd_sc_hd__a2bb2o_1
X_5953_ _1831_ _1876_ _1875_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__a21o_1
X_4904_ _0791_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5884_ _1760_ _1808_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__and2_1
X_8672_ net111 _3616_ vssd1 vssd1 vccd1 vccd1 _4123_ sky130_fd_sc_hd__xor2_1
X_4835_ _0709_ net87 vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__nand2_2
XFILLER_0_29_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7623_ allocation.game.lcdOutput.framebufferIndex\[12\] allocation.game.lcdOutput.framebufferIndex\[13\]
+ net120 vssd1 vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9283__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4766_ net89 _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__or2_1
X_7554_ net337 allocation.game.lcdOutput.tft.spi.data\[1\] net256 vssd1 vssd1 vccd1
+ vccd1 _0242_ sky130_fd_sc_hd__mux2_1
X_6505_ _0609_ _0610_ _2413_ net238 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4697_ net219 _0618_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7485_ _3058_ _3092_ _3099_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__a21oi_1
X_6436_ _2333_ _2348_ _2358_ _2343_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__o31a_1
X_9224_ clknet_leaf_22_clk _0037_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_9155_ clknet_leaf_12_clk _0217_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.color\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_6367_ allocation.game.cactusHeight1\[4\] allocation.game.cactusHeight1\[3\] _2279_
+ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5318_ _1174_ _1190_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__or2_1
X_8106_ _0613_ _2374_ vssd1 vssd1 vccd1 vccd1 _3608_ sky130_fd_sc_hd__and2_1
XANTENNA__4894__A1 _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9086_ clknet_leaf_14_clk _0182_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold13 _0244_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd3_1
X_6298_ allocation.game.controller.drawBlock.counter\[14\] _2180_ _2222_ vssd1 vssd1
+ vccd1 vccd1 _2223_ sky130_fd_sc_hd__a21bo_1
Xhold46 allocation.game.controller.init_module.idx\[4\] vssd1 vssd1 vccd1 vccd1 net369
+ sky130_fd_sc_hd__dlygate4sd3_1
X_8037_ _3543_ _3545_ vssd1 vssd1 vccd1 vccd1 _3546_ sky130_fd_sc_hd__nand2_1
X_5249_ net82 _1126_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__xor2_2
Xhold24 _0246_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 allocation.game.cactus2size.clock_div_inst0.counter\[13\] vssd1 vssd1 vccd1
+ vccd1 net358 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold68 allocation.game.controller.drawBlock.init_done vssd1 vssd1 vccd1 vccd1 net391
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 allocation.game.lcdOutput.tft.spi.tft_sdi vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold79 allocation.game.cactus2size.clock_div_inst0.counter\[0\] vssd1 vssd1 vccd1
+ vccd1 net402 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_27_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8939_ net131 _2282_ _3312_ _4387_ vssd1 vssd1 vccd1 vccd1 _4388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7899__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5066__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9156__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload4_A clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8543__C net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4620_ allocation.game.controller.drawBlock.x_start\[5\] allocation.game.controller.drawBlock.x_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__and2b_1
XANTENNA__4799__B net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4551_ net273 allocation.game.controller.v\[3\] vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7270_ _2935_ _2936_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4482_ allocation.game.game.score\[6\] vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6221_ _0993_ _1033_ _1035_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8067__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6152_ _2061_ _2062_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__xor2_1
X_5103_ net72 _0746_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__or2_1
X_6083_ _2007_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__inv_2
X_5034_ _0821_ _0868_ _0841_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a21o_1
X_6985_ allocation.game.scoreCounter.clock_div.counter\[20\] _2725_ net92 vssd1 vssd1
+ vccd1 vccd1 _2727_ sky130_fd_sc_hd__o21ai_1
X_5936_ _1816_ _1859_ _1860_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__and3_1
X_8724_ _4163_ _4174_ vssd1 vssd1 vccd1 vccd1 _4175_ sky130_fd_sc_hd__nor2_1
X_8655_ _0673_ net98 _4104_ _4105_ vssd1 vssd1 vccd1 vccd1 _4106_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5867_ _1790_ _1791_ _0896_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__a21o_1
X_7606_ net438 _2591_ _3014_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4818_ _0709_ _0742_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__nand2_2
X_8586_ net119 _4035_ _4036_ net97 _4034_ vssd1 vssd1 vccd1 vccd1 _4037_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5798_ _0738_ net86 vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9029__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4749_ _0649_ net104 vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__nand2_1
X_7537_ allocation.game.lcdOutput.tft.state\[0\] _3143_ _3145_ _3019_ vssd1 vssd1
+ vccd1 vccd1 _3146_ sky130_fd_sc_hd__a31o_1
X_7468_ net249 _3053_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__nand2_1
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_6419_ _2338_ _2341_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__or2_1
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
X_9207_ _0145_ _0404_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__7813__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7399_ net247 net245 vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__nand2_2
X_9138_ clknet_leaf_18_clk _0202_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_9069_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[15\] net190 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[15\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__7805__B2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout44_X net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8554__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6770_ allocation.game.cactus2size.clock_div_inst1.counter\[7\] allocation.game.cactus2size.clock_div_inst1.counter\[6\]
+ allocation.game.cactus2size.clock_div_inst1.counter\[9\] allocation.game.cactus2size.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5721_ _0897_ _1644_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8440_ _3318_ _3864_ vssd1 vssd1 vccd1 vccd1 _3893_ sky130_fd_sc_hd__or2_1
X_5652_ _1555_ _1557_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8371_ net140 _3578_ vssd1 vssd1 vccd1 vccd1 _3833_ sky130_fd_sc_hd__nand2_1
X_4603_ net269 _0472_ _0479_ net151 vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__o31a_1
X_5583_ _1506_ _1507_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__nor2_1
X_7322_ allocation.game.controller.init_module.delay_counter\[22\] allocation.game.controller.init_module.delay_counter\[21\]
+ _2967_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__nand3_1
XANTENNA__9321__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4534_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7253_ _4456_ allocation.game.dinoJump.next_dinoY\[0\] _2922_ _2923_ vssd1 vssd1
+ vccd1 vccd1 _2924_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4465_ net130 vssd1 vssd1 vccd1 vccd1 _4454_ sky130_fd_sc_hd__inv_2
X_7184_ allocation.game.dinoJump.count\[4\] _2870_ _0471_ vssd1 vssd1 vccd1 vccd1
+ _2872_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6204_ _2125_ _2126_ _1330_ _1378_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__a211o_1
XANTENNA__9471__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6135_ _2056_ _2057_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__xor2_1
X_6066_ _1948_ _1950_ _1949_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__a21o_1
X_5017_ _0940_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__or2_1
X_6968_ _2715_ _2716_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__nor2_1
X_8707_ _4151_ _4157_ vssd1 vssd1 vccd1 vccd1 _4158_ sky130_fd_sc_hd__or2_1
XANTENNA__7808__B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4785__B1 _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6899_ allocation.game.cactusDist.clock_div_inst0.counter\[0\] net155 _2673_ vssd1
+ vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__and3b_1
XANTENNA__8515__A2 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5919_ _1795_ _1842_ _1841_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8638_ _4083_ _4085_ _4088_ vssd1 vssd1 vccd1 vccd1 _4089_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8569_ _3298_ _4019_ _4016_ vssd1 vssd1 vccd1 vccd1 _4020_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9344__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9494__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7940_ allocation.game.controller.init_module.idx\[0\] _0425_ _2825_ _0398_ vssd1
+ vssd1 vccd1 vccd1 _3459_ sky130_fd_sc_hd__a31o_1
X_7871_ allocation.game.controller.drawBlock.counter\[1\] net108 net94 _3411_ vssd1
+ vssd1 vccd1 vccd1 _3412_ sky130_fd_sc_hd__a22o_1
X_6822_ allocation.game.cactus2size.clock_div_inst0.counter\[3\] _2622_ vssd1 vssd1
+ vccd1 vccd1 _2623_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6753_ allocation.game.cactus1size.clock_div_inst0.counter\[7\] allocation.game.cactus1size.clock_div_inst0.counter\[8\]
+ _2573_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__and3_1
X_9472_ clknet_leaf_12_clk _0379_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_end\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5704_ _1628_ _1627_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6684_ allocation.game.cactus1size.clock_div_inst1.counter\[1\] allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5635_ _1559_ _1552_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__nand2b_1
X_8423_ _3345_ net70 _3873_ vssd1 vssd1 vccd1 vccd1 _3876_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_21_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 allocation.game.controller.color\[10\] vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__dlygate4sd3_1
X_8354_ _0484_ _0509_ _3815_ _3816_ net136 vssd1 vssd1 vccd1 vccd1 _3817_ sky130_fd_sc_hd__o311a_1
XFILLER_0_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5566_ _1449_ _1450_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7305_ allocation.game.controller.init_module.delay_counter\[16\] allocation.game.controller.init_module.delay_counter\[15\]
+ _2956_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__and3_1
Xhold132 allocation.game.dinoJump.count\[19\] vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__dlygate4sd3_1
X_8285_ _2282_ net100 vssd1 vssd1 vccd1 vccd1 _3752_ sky130_fd_sc_hd__nor2_1
Xhold143 allocation.game.cactus1size.clock_div_inst0.counter\[12\] vssd1 vssd1 vccd1
+ vccd1 net466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 allocation.game.dinoJump.dinoDelay\[5\] vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4517_ allocation.game.dinoJump.dinoDelay\[3\] allocation.game.dinoJump.dinoDelay\[2\]
+ allocation.game.dinoJump.dinoDelay\[4\] allocation.game.dinoJump.dinoDelay\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__or4b_1
X_5497_ _1417_ _1420_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7236_ allocation.game.dinoJump.count\[15\] _2884_ _2899_ _2908_ vssd1 vssd1 vccd1
+ vccd1 _2909_ sky130_fd_sc_hd__and4_1
Xhold154 allocation.game.controller.init_module.delay_counter\[5\] vssd1 vssd1 vccd1
+ vccd1 net477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7167_ _2861_ _2862_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7098_ allocation.game.controller.drawBlock.y_start\[6\] _2787_ vssd1 vssd1 vccd1
+ vccd1 _2812_ sky130_fd_sc_hd__and2_1
X_6118_ _1957_ _1995_ _1996_ _1998_ _1985_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__a32o_1
XANTENNA__9217__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6049_ _1932_ _1933_ _1927_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__a21bo_1
XANTENNA__9367__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5521__B _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7729__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5249__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5420_ _0834_ _1198_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__nand2_1
X_5351_ _1274_ _1275_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8070_ _3502_ _3568_ _3577_ net204 net418 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__o32a_1
X_5282_ _1206_ _0917_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7021_ _0446_ _2750_ allocation.game.scoreCounter.bcd_tens\[1\] vssd1 vssd1 vccd1
+ vccd1 net19 sky130_fd_sc_hd__a21o_1
X_8972_ _2240_ net41 vssd1 vssd1 vccd1 vccd1 _4421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7923_ net95 _3446_ _3448_ net109 allocation.game.controller.drawBlock.counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7854_ _2778_ _2785_ allocation.game.controller.drawBlock.state\[2\] vssd1 vssd1
+ vccd1 vccd1 _3401_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7785_ _3308_ _3318_ vssd1 vssd1 vccd1 vccd1 _3347_ sky130_fd_sc_hd__nor2_1
X_6805_ allocation.game.cactus2size.clock_div_inst1.counter\[12\] _2610_ vssd1 vssd1
+ vccd1 vccd1 _2611_ sky130_fd_sc_hd__and2_1
X_4997_ _0798_ _0921_ _0893_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__a21o_1
X_9524_ net309 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_6736_ allocation.game.cactus1size.clock_div_inst0.counter\[1\] allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ allocation.game.cactus1size.clock_div_inst0.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2566_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6667_ _0620_ _2519_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9455_ clknet_leaf_18_clk _0362_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_8406_ allocation.game.controller.v\[7\] _3857_ vssd1 vssd1 vccd1 vccd1 _3860_ sky130_fd_sc_hd__xor2_1
X_9386_ clknet_leaf_13_clk _0296_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.idx\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_6598_ _2475_ _2476_ _2462_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[8\]
+ sky130_fd_sc_hd__and3b_1
X_5618_ _0810_ _1536_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__xor2_1
X_8337_ _0486_ _3799_ net139 vssd1 vssd1 vccd1 vccd1 _3801_ sky130_fd_sc_hd__a21oi_1
X_5549_ _1468_ _1471_ _1472_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8268_ net234 _3736_ net233 vssd1 vssd1 vccd1 vccd1 _3739_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9403__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7219_ _0471_ _2895_ _2897_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__and3_1
X_8199_ _0680_ _3688_ _0683_ vssd1 vssd1 vccd1 vccd1 _3689_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7393__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout71 _0801_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_4
Xfanout60 _0925_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_4
Xfanout82 net83 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8342__B1 allocation.game.controller.drawBlock.y_end\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout93 _2404_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_1
XFILLER_0_25_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8827__B _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7731__B net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9004__A _0462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _0842_ _0844_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4851_ _0572_ _0574_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_47_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_14_clk_X clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4782_ _0705_ _0706_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__and2b_4
X_7570_ net380 _3157_ _2526_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6521_ net444 _2421_ _2415_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__o21ai_1
X_6452_ _2344_ _2371_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9240_ clknet_leaf_22_clk _0024_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9171_ clknet_leaf_15_clk net53 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spiDataSet
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9062__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5403_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__inv_2
X_8122_ net239 _0615_ _3622_ _3597_ vssd1 vssd1 vccd1 vccd1 _3623_ sky130_fd_sc_hd__a31o_1
X_6383_ _2301_ _2298_ _2297_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__and3b_1
X_5334_ _1030_ _1237_ _1239_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__a21oi_1
X_8053_ _4459_ _3539_ vssd1 vssd1 vccd1 vccd1 _3561_ sky130_fd_sc_hd__nand2_1
X_5265_ _1181_ _1188_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__xnor2_1
X_5196_ _0733_ _1120_ _0725_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__o21a_1
X_7004_ _2739_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8955_ _3248_ _3256_ _4403_ _4026_ vssd1 vssd1 vccd1 vccd1 _4404_ sky130_fd_sc_hd__or4b_1
X_7906_ net95 _3435_ _3436_ net109 allocation.game.controller.drawBlock.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__a32o_1
X_8886_ _4262_ _4266_ _4335_ _4272_ vssd1 vssd1 vccd1 vccd1 _4336_ sky130_fd_sc_hd__a31o_1
X_7837_ net244 net242 net237 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7768_ _3301_ _3329_ _3323_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9507_ net292 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
X_7699_ _3251_ _3259_ _3254_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__o21bai_1
XANTENNA__9405__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6719_ net158 _2552_ _2553_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__nor3_1
Xclkload2 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9438_ clknet_leaf_12_clk _0347_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_9502__287 vssd1 vssd1 vccd1 vccd1 _9502__287/HI net287 sky130_fd_sc_hd__conb_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9369_ clknet_leaf_5_clk _0018_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.bcd_tens\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5352__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 allocation.game.lcdOutput.tft.initSeqCounter\[3\] vssd1 vssd1 vccd1 vccd1
+ net250 sky130_fd_sc_hd__clkbuf_2
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 allocation.game.collision.dinoY\[3\] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout74_X net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9085__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6630__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9325__RESET_B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8838__A net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5050_ _0780_ _0838_ _0940_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7189__A _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5952_ _1831_ _1875_ _1876_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__nand3_1
XANTENNA__6093__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8740_ net69 _4188_ _4190_ _3200_ vssd1 vssd1 vccd1 vccd1 _4191_ sky130_fd_sc_hd__o22a_1
X_4903_ _0826_ _0827_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__and2_1
XANTENNA__9428__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5883_ _0912_ _1645_ _1759_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__nand3_1
X_8671_ _0641_ _3616_ vssd1 vssd1 vccd1 vccd1 _4122_ sky130_fd_sc_hd__nand2_1
X_4834_ _0756_ _0757_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__xor2_2
X_7622_ _3183_ vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4765_ net105 _0691_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__or2_1
X_7553_ net331 allocation.game.lcdOutput.tft.spi.data\[0\] net256 vssd1 vssd1 vccd1
+ vccd1 _0241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6504_ net244 net163 vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8306__B1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout219_A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4696_ net219 net218 _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__or3_1
X_9223_ clknet_leaf_22_clk _0036_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_7484_ _3060_ _3095_ _3097_ _3098_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__a211o_1
X_6435_ _2353_ _2356_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6366_ _2285_ _2289_ _2288_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__or3b_1
X_9154_ clknet_leaf_3_clk _0216_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.clk1
+ sky130_fd_sc_hd__dfxtp_1
X_9085_ clknet_leaf_14_clk _0181_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5317_ _1232_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__nor2_1
XANTENNA__4894__A2 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8105_ _0688_ _3606_ vssd1 vssd1 vccd1 vccd1 _3607_ sky130_fd_sc_hd__or2_1
X_8036_ _3544_ vssd1 vssd1 vccd1 vccd1 _3545_ sky130_fd_sc_hd__inv_2
Xhold14 allocation.game.lcdOutput.tft.spi.dataShift\[6\] vssd1 vssd1 vccd1 vccd1 net337
+ sky130_fd_sc_hd__dlygate4sd3_1
X_6297_ allocation.game.controller.drawBlock.counter\[14\] _2180_ _2181_ allocation.game.controller.drawBlock.counter\[13\]
+ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__o221a_1
Xhold47 allocation.game.controller.init_module.idx\[5\] vssd1 vssd1 vccd1 vccd1 net370
+ sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _1171_ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__and2b_1
Xhold36 allocation.game.lcdOutput.tft.spi.data\[6\] vssd1 vssd1 vccd1 vccd1 net359
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 allocation.game.dinoJump.dinoDelay\[20\] vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _0930_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__nor2_1
Xhold69 _0293_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 allocation.game.scoreCounter.clock_div.counter\[1\] vssd1 vssd1 vccd1 vccd1
+ net381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5900__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8938_ net133 _4386_ _2278_ vssd1 vssd1 vccd1 vccd1 _4387_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_27_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8869_ _4318_ vssd1 vssd1 vccd1 vccd1 _4319_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4885__A2 _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7737__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5257__A _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4550_ net273 allocation.game.controller.v\[3\] vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4481_ allocation.game.game.score\[1\] vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__inv_2
X_6220_ _2143_ _2144_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8067__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6151_ _2075_ _2074_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__and2b_1
XANTENNA__9100__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5102_ net72 _0746_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6082_ _1969_ _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__nand3_1
X_5033_ _0956_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__nand2_1
XANTENNA__9250__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6984_ _2725_ _2726_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout169_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5935_ _1813_ _1815_ _1814_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__a21o_1
X_8723_ net142 net57 _4173_ vssd1 vssd1 vccd1 vccd1 _4174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8654_ net89 net116 vssd1 vssd1 vccd1 vccd1 _4105_ sky130_fd_sc_hd__nor2_1
X_5866_ _1740_ _1789_ _1788_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__a21o_1
X_4817_ _0741_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7605_ net143 _3175_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8585_ net217 _4031_ vssd1 vssd1 vccd1 vccd1 _4036_ sky130_fd_sc_hd__nand2_1
X_5797_ _1670_ _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4748_ net89 net104 vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__nand2_2
X_7536_ _0429_ net252 _3144_ net245 vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_47_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4679_ net2 net1 net5 vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nand3b_1
X_7467_ _4463_ net252 vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__nand2_2
X_6418_ _0422_ allocation.game.game.score\[5\] allocation.game.scoreCounter.clock_div.slow_clk
+ _2324_ _2340_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__o41a_1
X_9206_ _0144_ _0403_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__7813__C net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__clkbuf_4
X_9137_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[31\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[31\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7398_ allocation.game.lcdOutput.tft.state\[0\] _3018_ vssd1 vssd1 vccd1 vccd1 _3020_
+ sky130_fd_sc_hd__nand2_2
X_6349_ net164 _0654_ _0652_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__o21a_1
X_9068_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[14\] net190 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[14\] sky130_fd_sc_hd__dfrtp_1
X_8019_ _0491_ _0499_ vssd1 vssd1 vccd1 vccd1 _3529_ sky130_fd_sc_hd__nor2_1
XANTENNA__5630__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout37_X net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8005__X _3516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9508__293 vssd1 vssd1 vccd1 vccd1 _9508__293/HI net293 sky130_fd_sc_hd__conb_1
XANTENNA__4533__X _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8297__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9123__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9273__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9012__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5720_ _0896_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5651_ _1533_ _1561_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__xnor2_1
X_8370_ _0541_ _3580_ _3816_ net139 vssd1 vssd1 vccd1 vccd1 _3832_ sky130_fd_sc_hd__a31o_1
X_4602_ _0534_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoY\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_26_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5582_ _1492_ _1504_ _1505_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__nor3_1
X_7321_ allocation.game.controller.init_module.delay_counter\[21\] _2967_ allocation.game.controller.init_module.delay_counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__a21o_1
XANTENNA__8298__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4533_ _0465_ _0470_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__or2_4
X_7252_ _4456_ allocation.game.dinoJump.next_dinoY\[0\] _0538_ net268 _2918_ vssd1
+ vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_29_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4464_ allocation.game.lcdOutput.framebufferIndex\[0\] vssd1 vssd1 vccd1 vccd1 _0401_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6203_ _1378_ _2127_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__nor2_1
X_7183_ _0472_ _2870_ _2871_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__nor3_1
XFILLER_0_42_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6134_ net103 _0895_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__nor2_1
X_6065_ _1987_ _1988_ _1986_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__a21bo_1
X_5016_ _0802_ _0939_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6967_ net467 _2713_ net93 vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__o21ai_1
X_8706_ net111 _3670_ vssd1 vssd1 vccd1 vccd1 _4157_ sky130_fd_sc_hd__and2_1
X_5918_ _1795_ _1841_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6898_ _2673_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__inv_2
X_8637_ net99 _4084_ _4086_ _4087_ vssd1 vssd1 vccd1 vccd1 _4088_ sky130_fd_sc_hd__o31a_1
X_5849_ _1767_ _1773_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__nor2_1
XANTENNA__9146__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8568_ _4017_ _4018_ _0611_ vssd1 vssd1 vccd1 vccd1 _4019_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7519_ net345 _3130_ net53 vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8499_ net126 _3311_ _3950_ _3271_ vssd1 vssd1 vccd1 vccd1 _3951_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9296__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7840__A _2973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7839__X _3394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8978__B1 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7870_ allocation.game.controller.drawBlock.counter\[0\] allocation.game.controller.drawBlock.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3411_ sky130_fd_sc_hd__nand2_1
X_6821_ net161 _2621_ _2622_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_34_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_15_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
X_6752_ allocation.game.cactus1size.clock_div_inst0.counter\[7\] _2573_ allocation.game.cactus1size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__a21oi_1
X_9471_ clknet_leaf_11_clk _0378_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_end\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_5703_ _0750_ _1620_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__xor2_1
X_6683_ allocation.game.det allocation.game.dinoJump.button vssd1 vssd1 vccd1 vccd1
+ _2529_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5634_ _1553_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__xnor2_1
X_8422_ _3345_ net70 _3873_ vssd1 vssd1 vccd1 vccd1 _3875_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_21_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8353_ _0484_ _3815_ _0509_ vssd1 vssd1 vccd1 vccd1 _3816_ sky130_fd_sc_hd__o21ai_1
X_7304_ net428 _2956_ _2958_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__o21a_1
Xhold100 _0104_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__dlygate4sd3_1
X_5565_ _1487_ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold144 allocation.game.scoreCounter.clock_div.counter\[13\] vssd1 vssd1 vccd1 vccd1
+ net467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold111 allocation.game.controller.drawBlock.x_end\[3\] vssd1 vssd1 vccd1 vccd1 net434
+ sky130_fd_sc_hd__dlygate4sd3_1
X_8284_ net81 _2256_ vssd1 vssd1 vccd1 vccd1 _3751_ sky130_fd_sc_hd__nor2_1
Xhold133 allocation.game.cactusDist.clock_div_inst0.counter\[6\] vssd1 vssd1 vccd1
+ vccd1 net456 sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ allocation.game.dinoJump.dinoDelay\[1\] allocation.game.dinoJump.dinoDelay\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__or2_1
Xhold122 allocation.game.cactus2size.clock_div_inst1.counter\[12\] vssd1 vssd1 vccd1
+ vccd1 net445 sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ net61 _1374_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__xnor2_1
X_7235_ allocation.game.dinoJump.count\[16\] allocation.game.dinoJump.count\[17\]
+ allocation.game.dinoJump.count\[18\] vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_1_0__f_clk_X clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold155 allocation.game.cactusDist.clock_div_inst1.counter\[6\] vssd1 vssd1 vccd1
+ vccd1 net478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7166_ _0401_ net132 vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__or2_1
X_6117_ _2040_ _2041_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__and2b_1
X_7097_ _2802_ _2809_ _2811_ _2801_ vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__o31a_1
X_6048_ _1970_ _1972_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7999_ net274 _3487_ _3509_ net137 vssd1 vssd1 vccd1 vccd1 _3510_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4997__A1 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9311__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9461__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8360__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5350_ _1270_ _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand3_1
X_5281_ _0797_ _0921_ _1205_ _0893_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7020_ allocation.game.scoreCounter.bcd_tens\[2\] _2748_ _2749_ vssd1 vssd1 vccd1
+ vccd1 _2750_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_4_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
X_9530__312 vssd1 vssd1 vccd1 vccd1 _9530__312/HI net312 sky130_fd_sc_hd__conb_1
X_8971_ _2249_ net45 _4419_ vssd1 vssd1 vccd1 vccd1 _4420_ sky130_fd_sc_hd__o21ai_1
X_7922_ _3447_ vssd1 vssd1 vccd1 vccd1 _3448_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7853_ allocation.game.controller.drawBlock.idx\[3\] allocation.game.controller.drawBlock.idx\[2\]
+ _2769_ allocation.game.controller.drawBlock.idx\[4\] vssd1 vssd1 vccd1 vccd1 _3400_
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__7639__B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7926__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout151_A _0462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4996_ _0920_ _0889_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__and2b_1
X_6804_ net158 _2609_ _2610_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__nor3_1
X_7784_ net118 _3296_ _3345_ _3344_ vssd1 vssd1 vccd1 vccd1 _3346_ sky130_fd_sc_hd__o31a_1
X_9523_ net308 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
X_6735_ allocation.game.cactus1size.clock_div_inst0.counter\[1\] allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ allocation.game.cactus1size.clock_div_inst0.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2565_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9454_ clknet_leaf_18_clk _0361_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_6666_ net229 net228 allocation.game.cactusMove.pixel\[4\] vssd1 vssd1 vccd1 vccd1
+ _2519_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8405_ allocation.game.controller.v\[7\] net85 vssd1 vssd1 vccd1 vccd1 _3859_ sky130_fd_sc_hd__nand2_1
X_6597_ allocation.game.cactusMove.count\[7\] _2472_ allocation.game.cactusMove.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__a21o_1
X_9385_ clknet_leaf_13_clk _0295_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.idx\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5617_ _0777_ _0892_ _1540_ _1538_ _1494_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8336_ _0486_ _3799_ vssd1 vssd1 vccd1 vccd1 _3800_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5548_ _1468_ _1471_ _1472_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8267_ net145 net153 _3737_ vssd1 vssd1 vccd1 vccd1 _3738_ sky130_fd_sc_hd__a21oi_1
X_7218_ _2896_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__inv_2
X_5479_ _1385_ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__xnor2_1
X_8198_ _0663_ _0678_ vssd1 vssd1 vccd1 vccd1 _3688_ sky130_fd_sc_hd__or2_1
X_7149_ _2841_ _2851_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__nand2_1
XANTENNA__9334__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7614__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout64_A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9484__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout72 _0726_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_4
Xfanout83 _0714_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_2
Xfanout50 _3228_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_4
Xfanout61 net62 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout94 net95 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_2
XFILLER_0_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9004__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7081__A1 allocation.game.controller.drawBlock.y_end\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9020__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4850_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_0_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4781_ _0579_ _0601_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_32_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6520_ allocation.game.dinoJump.dinoDelay\[4\] allocation.game.dinoJump.dinoDelay\[5\]
+ _2419_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4611__B _0541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6451_ _2348_ _2363_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__nor2_1
X_6382_ net274 _2280_ _2305_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__a21oi_1
X_9170_ clknet_leaf_15_clk _0232_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_5402_ _1323_ _1325_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__nand3_2
X_8121_ net224 _0612_ vssd1 vssd1 vccd1 vccd1 _3622_ sky130_fd_sc_hd__nand2_1
X_5333_ _1207_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9357__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8052_ _4459_ _3539_ vssd1 vssd1 vccd1 vccd1 _3560_ sky130_fd_sc_hd__or2_2
X_5264_ _1188_ _1181_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nand2b_1
X_5195_ _0727_ _0761_ _0782_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__a21oi_1
X_7003_ _0451_ _2737_ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8954_ _4027_ _4080_ _4399_ _4402_ vssd1 vssd1 vccd1 vccd1 _4403_ sky130_fd_sc_hd__or4b_1
X_7905_ allocation.game.controller.drawBlock.counter\[9\] allocation.game.controller.drawBlock.counter\[10\]
+ _3427_ allocation.game.controller.drawBlock.counter\[11\] vssd1 vssd1 vccd1 vccd1
+ _3436_ sky130_fd_sc_hd__a31o_1
X_8885_ _4300_ _4229_ vssd1 vssd1 vccd1 vccd1 _4335_ sky130_fd_sc_hd__and2b_1
X_7836_ net461 allocation.game.controller.state\[0\] net237 vssd1 vssd1 vccd1 vccd1
+ _0285_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4979_ _0700_ _0902_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__or2_2
X_7767_ _3299_ _3308_ _3326_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__or3_1
X_9506_ net291 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XANTENNA__8324__A1 _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4802__A _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_4
X_7698_ _3251_ _3259_ _3254_ vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__o21ba_1
X_6718_ allocation.game.cactus1size.clock_div_inst1.counter\[11\] allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ _2549_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9437_ clknet_leaf_12_clk _0346_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__9373__Q allocation.game.controller.drawBlock.state\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6649_ _2507_ _2508_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[27\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9368_ clknet_leaf_5_clk _0017_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.bcd_tens\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_8319_ _3782_ _3783_ net134 vssd1 vssd1 vccd1 vccd1 _3784_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9299_ clknet_leaf_22_clk _0085_ net180 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout240 allocation.game.controller.state\[9\] vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout273 allocation.game.collision.dinoY\[3\] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout251 allocation.game.lcdOutput.tft.initSeqCounter\[2\] vssd1 vssd1 vccd1 vccd1
+ net251 sky130_fd_sc_hd__buf_2
XANTENNA_fanout67_X net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4585__C1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7669__A3 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9015__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8854__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5951_ _1828_ _1830_ _1829_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4902_ _0818_ _0825_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8670_ _4091_ _4119_ _4120_ net46 vssd1 vssd1 vccd1 vccd1 _4121_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5882_ _1803_ _1806_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4833_ _0756_ _0757_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__and2_4
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7621_ allocation.game.lcdOutput.framebufferIndex\[12\] net120 vssd1 vssd1 vccd1
+ vccd1 _3183_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4764_ net112 _0658_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7552_ net247 _3043_ _3149_ net245 vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__a31o_1
X_6503_ allocation.game.controller.state\[6\] allocation.game.controller.state\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__or2_1
X_7483_ net247 net245 _3048_ _3020_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4695_ net222 _0621_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6434_ _2356_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9222_ clknet_leaf_22_clk _0035_ net169 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout114_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9153_ clknet_leaf_13_clk _0400_ net210 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6365_ _4457_ _2278_ _2286_ _0436_ _4456_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9084_ clknet_leaf_14_clk _0180_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_5316_ _1239_ _1240_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__or2_1
X_8104_ net142 _0686_ vssd1 vssd1 vccd1 vccd1 _3606_ sky130_fd_sc_hd__and2_1
X_6296_ allocation.game.controller.drawBlock.counter\[12\] _2183_ _2220_ _2182_ vssd1
+ vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__o211a_1
X_8035_ allocation.game.controller.v\[5\] _3541_ vssd1 vssd1 vccd1 vccd1 _3544_ sky130_fd_sc_hd__and2_1
X_5247_ _1169_ _1170_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__or2_1
Xhold37 allocation.game.lcdOutput.tft.spi.dataDc vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 allocation.game.cactusMove.count\[31\] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 _0242_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5178_ _0884_ _0929_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__and2_1
Xhold59 _0116_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold48 allocation.game.lcdOutput.tft.remainingDelayTicks\[9\] vssd1 vssd1 vccd1 vccd1
+ net371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8937_ _0401_ allocation.game.cactusHeight1\[0\] allocation.game.cactusHeight1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _4386_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_27_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8868_ _4316_ _4317_ vssd1 vssd1 vccd1 vccd1 _4318_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_17_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5359__A1 _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7819_ _2353_ _2372_ vssd1 vssd1 vccd1 vccd1 _3378_ sky130_fd_sc_hd__nor2_1
X_8799_ _4229_ _4248_ _4246_ vssd1 vssd1 vccd1 vccd1 _4249_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5628__A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7562__B _2526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8674__A _0673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_X clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9052__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7737__B net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7753__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4480_ allocation.game.lcdOutput.tft.state\[0\] vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6150_ _2059_ _2060_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5101_ _0830_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6081_ _1967_ _1968_ _0712_ _0729_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__a2bb2o_1
X_5032_ _0875_ _0877_ _0955_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__nand3_1
X_6983_ allocation.game.scoreCounter.clock_div.counter\[19\] _2724_ net92 vssd1 vssd1
+ vccd1 vccd1 _2726_ sky130_fd_sc_hd__o21ai_1
X_5934_ _0716_ _0885_ _1858_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__and3_1
X_8722_ _0657_ _3228_ _3668_ net57 vssd1 vssd1 vccd1 vccd1 _4173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8653_ _0669_ _0670_ net116 vssd1 vssd1 vccd1 vccd1 _4104_ sky130_fd_sc_hd__and3_1
X_5865_ _1740_ _1788_ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__nand3_1
X_4816_ _0720_ _0734_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7604_ allocation.game.cactusDist.lfsr2\[1\] allocation.game.cactusDist.lfsr2\[0\]
+ allocation.game.cactusDist.clock_div_inst1.clk1 vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8584_ net217 _4031_ vssd1 vssd1 vccd1 vccd1 _4035_ sky130_fd_sc_hd__or2_1
X_5796_ net110 _0887_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7535_ _3093_ _3119_ _3131_ net247 vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4747_ _0669_ _0670_ net104 vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__and3_1
X_4678_ _0417_ allocation.game.controller.drawBlock.state\[2\] _0606_ _0607_ vssd1
+ vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a22o_1
X_7466_ net250 _3052_ vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6417_ _2336_ _2339_ allocation.game.game.score\[6\] vssd1 vssd1 vccd1 vccd1 _2340_
+ sky130_fd_sc_hd__a21o_1
X_9205_ _0143_ _0402_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_7397_ allocation.game.lcdOutput.tft.state\[2\] allocation.game.lcdOutput.tft.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__nand2b_2
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6348_ _2252_ _2270_ _2271_ _2269_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__a31o_1
X_9136_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[30\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[30\] sky130_fd_sc_hd__dfrtp_1
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9067_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[13\] net192 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[13\] sky130_fd_sc_hd__dfrtp_1
X_6279_ _2092_ _2203_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__or2_1
X_8018_ _3494_ _3527_ vssd1 vssd1 vccd1 vccd1 _3528_ sky130_fd_sc_hd__nor2_1
XANTENNA__9075__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5504__A1 _0729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9418__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8757__A1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_5650_ _1574_ _1573_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__and2b_1
X_4601_ net273 _0481_ _0533_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5581_ _1492_ _1504_ _1505_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__o21a_1
X_7320_ allocation.game.controller.init_module.delay_counter\[21\] _2967_ _2968_ vssd1
+ vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__o21a_1
X_4532_ _4456_ net258 _0468_ _0469_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or4_2
XANTENNA__9471__Q allocation.game.controller.drawBlock.y_end\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7251_ net269 _0538_ _2920_ _2921_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6202_ _2125_ _2126_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__and2_1
XANTENNA__9098__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7182_ net148 _2868_ allocation.game.dinoJump.count\[3\] vssd1 vssd1 vccd1 vccd1
+ _2871_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6133_ _2056_ _2057_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__and2_1
XANTENNA_clkload16_A clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6064_ _1986_ _1988_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__nand2_1
X_5015_ _0802_ _0939_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout181_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6966_ allocation.game.scoreCounter.clock_div.counter\[13\] allocation.game.scoreCounter.clock_div.counter\[12\]
+ _2712_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5917_ _1792_ _1793_ _1794_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8705_ net120 _4154_ _4155_ net98 vssd1 vssd1 vccd1 vccd1 _4156_ sky130_fd_sc_hd__a22o_1
XANTENNA__4785__A2 _0708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6897_ _2670_ _2672_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7184__B1 _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8636_ _3999_ _4086_ net99 vssd1 vssd1 vccd1 vccd1 _4087_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8920__A1 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5848_ _1769_ _1772_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5779_ net82 _1596_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__and2b_1
X_8567_ net227 net52 vssd1 vssd1 vccd1 vccd1 _4018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7518_ _3110_ _3128_ _3129_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8498_ net130 _0442_ _3311_ _3312_ vssd1 vssd1 vccd1 vccd1 _3950_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7449_ allocation.game.lcdOutput.r_over allocation.game.lcdOutput.r_idle allocation.game.lcdOutput.r_win
+ allocation.game.lcdOutput.r_cloud vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__or4_2
XANTENNA__8936__B net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout94_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9119_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[13\] net173 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__7840__B _3394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6737__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8952__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9240__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9023__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9390__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5551__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9524__309 vssd1 vssd1 vccd1 vccd1 _9524__309/HI net309 sky130_fd_sc_hd__conb_1
X_6820_ allocation.game.cactus2size.clock_div_inst0.counter\[0\] allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ allocation.game.cactus2size.clock_div_inst0.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2622_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_19_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6751_ allocation.game.cactus1size.clock_div_inst0.counter\[7\] _2573_ _2575_ vssd1
+ vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__o21a_1
XANTENNA__5964__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9470_ clknet_leaf_11_clk _0377_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_end\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5702_ net88 _0892_ _1626_ _1623_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__a31o_1
X_6682_ allocation.game.det allocation.game.dinoJump.button vssd1 vssd1 vccd1 vccd1
+ _2528_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5633_ _1555_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__and2_1
X_8421_ net119 _3872_ vssd1 vssd1 vccd1 vccd1 _3874_ sky130_fd_sc_hd__nand2_1
X_8352_ _0483_ _3799_ vssd1 vssd1 vccd1 vccd1 _3815_ sky130_fd_sc_hd__nor2_1
X_5564_ _1436_ _1488_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__nand2_1
X_7303_ net123 _2957_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__nor2_1
Xhold101 allocation.game.scoreCounter.clock_div.counter\[15\] vssd1 vssd1 vccd1 vccd1
+ net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4515_ _0452_ _0453_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8283_ allocation.game.controller.drawBlock.y_end\[1\] net196 _3749_ _3750_ vssd1
+ vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__o22a_1
Xhold134 allocation.game.cactusMove.count\[30\] vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 allocation.game.cactus1size.clock_div_inst0.counter\[4\] vssd1 vssd1 vccd1
+ vccd1 net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 allocation.game.cactus2size.clock_div_inst1.counter\[9\] vssd1 vssd1 vccd1
+ vccd1 net446 sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ net61 _1419_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__nand2_1
Xhold156 allocation.game.scoreCounter.clock_div.counter\[9\] vssd1 vssd1 vccd1 vccd1
+ net479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7234_ _4461_ _2906_ _2907_ net84 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold145 allocation.game.dinoJump.dinoDelay\[16\] vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7165_ _0401_ net132 vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__nand2_1
XANTENNA__8969__B2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6116_ _2012_ _2039_ _2038_ _2035_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__o211ai_1
X_7096_ allocation.game.controller.drawBlock.y_end\[5\] _2779_ _2787_ allocation.game.controller.drawBlock.y_start\[5\]
+ _2810_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__a221o_1
X_6047_ _1967_ _1970_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__nand3_1
XANTENNA__4805__A _0729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7388__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7998_ net274 _3487_ vssd1 vssd1 vccd1 vccd1 _3509_ sky130_fd_sc_hd__nor2_1
XANTENNA__9113__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6949_ allocation.game.scoreCounter.clock_div.counter\[7\] _2399_ vssd1 vssd1 vccd1
+ vccd1 _2704_ sky130_fd_sc_hd__nand2_1
XANTENNA__8354__C1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9263__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8619_ _0614_ _2375_ net75 vssd1 vssd1 vccd1 vccd1 _4070_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8409__B1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9319__RESET_B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7935__A2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6930__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9018__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8857__A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5280_ _0834_ _1201_ _1204_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8576__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8970_ net129 _2253_ net45 _2249_ _4418_ vssd1 vssd1 vccd1 vccd1 _4419_ sky130_fd_sc_hd__a221o_1
XANTENNA__9136__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7921_ allocation.game.controller.drawBlock.counter\[15\] allocation.game.controller.drawBlock.counter\[16\]
+ _3442_ vssd1 vssd1 vccd1 vccd1 _3447_ sky130_fd_sc_hd__and3_1
X_7852_ allocation.game.controller.block_done allocation.game.controller.drawBlock.state\[3\]
+ net236 vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ net86 _0919_ net79 vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9286__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6803_ allocation.game.cactus2size.clock_div_inst1.counter\[11\] allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ _2606_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__and3_1
X_7783_ net58 net51 vssd1 vssd1 vccd1 vccd1 _3345_ sky130_fd_sc_hd__nand2_1
X_9522_ net307 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6734_ net154 _2561_ _2563_ _2564_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__and4_1
X_9453_ clknet_leaf_18_clk _0360_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8404_ _3842_ _3858_ _3856_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__o21ai_1
X_6665_ net228 net226 vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9384_ clknet_leaf_13_clk _0294_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.block_done
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6596_ allocation.game.cactusMove.count\[7\] allocation.game.cactusMove.count\[8\]
+ _2472_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__and3_1
X_5616_ _1494_ _1538_ _1540_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__a21boi_1
X_8335_ _0503_ _3786_ vssd1 vssd1 vccd1 vccd1 _3799_ sky130_fd_sc_hd__and2_1
X_5547_ _1412_ _1414_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8266_ _2316_ _3735_ _3736_ net146 vssd1 vssd1 vccd1 vccd1 _3737_ sky130_fd_sc_hd__o211a_1
X_5478_ _1356_ _1402_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__and2_1
X_7217_ allocation.game.dinoJump.count\[13\] allocation.game.dinoJump.count\[12\]
+ _2891_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8197_ _3680_ _3682_ _3687_ net207 net410 vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__o32a_1
X_7148_ net125 _2840_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__or2_1
X_7079_ allocation.game.controller.drawBlock.idx\[4\] _2762_ _2771_ vssd1 vssd1 vccd1
+ vccd1 _2797_ sky130_fd_sc_hd__or3_1
XANTENNA__4806__Y _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout57_A _3219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 _3275_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_2
Xfanout73 _0726_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_1
XFILLER_0_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout62 net63 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_4
Xfanout51 _3227_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_12_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout84 _2863_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_2
XFILLER_0_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout95 _3410_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_2
XFILLER_0_9_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8677__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4780_ _0702_ _0703_ _0704_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__nand3_4
XANTENNA__6660__A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7756__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6450_ allocation.game.scoreCounter.bcd_tens\[2\] _2369_ _2370_ net147 vssd1 vssd1
+ vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
Xclkload10 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_12
XFILLER_0_3_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7541__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6381_ net274 _2280_ _2282_ net277 vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__o211a_1
X_5401_ net62 _1276_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__xnor2_1
X_8120_ _3620_ vssd1 vssd1 vccd1 vccd1 _3621_ sky130_fd_sc_hd__inv_2
X_5332_ _0917_ _1206_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8051_ _3501_ _3502_ _3559_ net203 net405 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__o32a_1
X_5263_ _1186_ _1187_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nand2_1
X_5194_ _1117_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__nand2b_1
X_7002_ _0450_ _0451_ _2738_ _2735_ _2734_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__o32a_1
X_8953_ _3208_ _3673_ _4400_ _4401_ vssd1 vssd1 vccd1 vccd1 _4402_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7904_ _3434_ vssd1 vssd1 vccd1 vccd1 _3435_ sky130_fd_sc_hd__inv_2
X_8884_ _4321_ _4331_ _4332_ _3873_ _4333_ vssd1 vssd1 vccd1 vccd1 _4334_ sky130_fd_sc_hd__o221a_1
X_7835_ net232 _3383_ _3392_ net234 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9505_ net290 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_4978_ _0700_ _0902_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7766_ net117 _3308_ vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload4 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload4/X sky130_fd_sc_hd__clkbuf_4
X_7697_ _3239_ _3258_ vssd1 vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__and2_1
X_6717_ allocation.game.cactus1size.clock_div_inst1.counter\[10\] _2549_ allocation.game.cactus1size.clock_div_inst1.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9436_ clknet_leaf_11_clk _0345_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6648_ allocation.game.cactusMove.count\[27\] _2506_ net150 vssd1 vssd1 vccd1 vccd1
+ _2508_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9367_ clknet_leaf_6_clk _0016_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.bcd_tens\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6579_ allocation.game.cactusMove.count\[1\] allocation.game.cactusMove.count\[0\]
+ allocation.game.cactusMove.count\[2\] vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__a21o_1
X_8318_ net273 _3761_ net268 vssd1 vssd1 vccd1 vccd1 _3783_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9301__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9298_ clknet_leaf_21_clk _0084_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_8249_ allocation.game.lcdOutput.tft.remainingDelayTicks\[13\] _2991_ allocation.game.lcdOutput.tft.remainingDelayTicks\[14\]
+ vssd1 vssd1 vccd1 vccd1 _3725_ sky130_fd_sc_hd__o21ai_1
Xfanout241 allocation.game.controller.state\[8\] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
Xfanout230 allocation.game.cactusMove.pixel\[2\] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5846__B1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout274 allocation.game.collision.dinoY\[3\] vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
Xfanout263 allocation.game.collision.dinoY\[6\] vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout252 allocation.game.lcdOutput.tft.initSeqCounter\[1\] vssd1 vssd1 vccd1 vccd1
+ net252 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5808__B _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6326__B2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5950_ _1871_ _1874_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__nand2_1
X_4901_ _0818_ _0825_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7620_ allocation.game.lcdOutput.framebufferIndex\[16\] _2843_ _3180_ vssd1 vssd1
+ vccd1 vccd1 _3182_ sky130_fd_sc_hd__o21ai_1
X_5881_ _1804_ _1805_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_16_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4832_ _0549_ _0570_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ net112 _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__and2_1
X_7551_ net247 _3153_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__xnor2_1
XANTENNA__9324__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6502_ allocation.game.controller.state\[6\] allocation.game.controller.state\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__nor2_2
X_4694_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__inv_2
X_7482_ _0429_ net245 _3084_ _3096_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__and4_1
X_6433_ _2318_ _2354_ _2355_ _2319_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__a2bb2o_2
X_9221_ clknet_leaf_22_clk _0047_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9152_ clknet_leaf_13_clk _0399_ net210 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout107_A _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6364_ net279 _2287_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9083_ clknet_leaf_14_clk _0179_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__9474__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8103_ _3597_ _3604_ _3605_ net203 net434 vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__o32a_1
X_5315_ _1236_ _1238_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__and2b_1
X_6295_ _2184_ _2186_ _2219_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8034_ allocation.game.controller.v\[5\] _3541_ vssd1 vssd1 vccd1 vccd1 _3543_ sky130_fd_sc_hd__or2_1
X_5246_ _1169_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__and2_1
Xhold38 allocation.game.lcdOutput.tft.spi.cs vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 allocation.game.lcdOutput.tft.spi.dataShift\[0\] vssd1 vssd1 vccd1 vccd1 net350
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 allocation.game.cactus1size.clock_div_inst1.counter\[13\] vssd1 vssd1 vccd1
+ vccd1 net339 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5177_ _1096_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__nor2_1
Xhold49 allocation.game.scoreCounter.clock_div.counter\[4\] vssd1 vssd1 vccd1 vccd1
+ net372 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8936_ _2294_ net37 vssd1 vssd1 vccd1 vccd1 _4385_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8867_ _4454_ net275 vssd1 vssd1 vccd1 vccd1 _4317_ sky130_fd_sc_hd__or2_1
X_7818_ allocation.game.bcd_ones\[1\] _2369_ _3377_ net146 vssd1 vssd1 vccd1 vccd1
+ _0282_ sky130_fd_sc_hd__a22o_1
X_8798_ net131 _3486_ _3760_ _4247_ vssd1 vssd1 vccd1 vccd1 _4248_ sky130_fd_sc_hd__a31o_1
XANTENNA__9384__Q allocation.game.controller.block_done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4532__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7749_ net42 net40 vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_7_Left_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9419_ clknet_leaf_11_clk _0328_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_start\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8955__A _3248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6492__B1 allocation.game.controller.drawBlock.state\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9347__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8270__A2_N net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8865__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5100_ _1023_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6080_ _2002_ _2004_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__nor2_1
X_5031_ _0875_ _0877_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9469__Q allocation.game.controller.drawBlock.y_end\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6982_ allocation.game.scoreCounter.clock_div.counter\[19\] _2724_ vssd1 vssd1 vccd1
+ vccd1 _2725_ sky130_fd_sc_hd__and2_1
X_8721_ _4165_ _4171_ vssd1 vssd1 vccd1 vccd1 _4172_ sky130_fd_sc_hd__nor2_1
X_5933_ net141 net86 vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_49_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8652_ _4102_ vssd1 vssd1 vccd1 vccd1 _4103_ sky130_fd_sc_hd__inv_2
X_5864_ _1738_ _1739_ _0901_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a21o_1
X_4815_ _0739_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__inv_2
X_8583_ _4031_ _4033_ vssd1 vssd1 vccd1 vccd1 _4034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7603_ _3173_ _3174_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5795_ net80 _1674_ _1719_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7534_ _0429_ _3142_ _3132_ net245 vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4746_ net104 vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4677_ allocation.game.controller.drawBlock.state\[0\] allocation.game.controller.drawBlock.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__or2_1
X_7465_ net249 _3076_ _3080_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6416_ allocation.game.game.score\[5\] allocation.game.game.score\[4\] _2330_ _0438_
+ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__a31o_1
X_9204_ _0142_ _0414_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_7396_ allocation.game.lcdOutput.tft.state\[2\] allocation.game.lcdOutput.tft.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__and2b_2
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__clkbuf_4
X_6347_ _2261_ _2262_ _2264_ _2259_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__and4b_1
X_9135_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[29\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8775__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5277__A1 _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9066_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[12\] net190 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[12\] sky130_fd_sc_hd__dfrtp_1
X_6278_ _2089_ _2091_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__nor2_1
X_8017_ _3503_ _3504_ vssd1 vssd1 vccd1 vccd1 _3527_ sky130_fd_sc_hd__nor2_1
X_5229_ net60 _1143_ _1146_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__nand3_1
XANTENNA__4527__B _0464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8919_ net41 _4353_ _4366_ net36 _4363_ vssd1 vssd1 vccd1 vccd1 _4369_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload2_A clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ net143 _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5580_ _1452_ _1453_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531_ net278 net268 _0466_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or3b_1
X_7250_ _4457_ allocation.game.dinoJump.next_dinoY\[1\] allocation.game.dinoJump.next_dinoY\[3\]
+ _4458_ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6201_ _1375_ _1377_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__xnor2_1
X_7181_ allocation.game.dinoJump.count\[3\] net148 _2868_ vssd1 vssd1 vccd1 vccd1
+ _2870_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6132_ _2023_ _2024_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__xor2_1
XANTENNA__8445__B2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6063_ _0712_ _0905_ _1946_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__a21o_1
XANTENNA__8996__A2 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5014_ _0780_ _0838_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout174_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6965_ _2713_ _2714_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__nor2_1
X_8704_ net104 _4151_ vssd1 vssd1 vccd1 vccd1 _4155_ sky130_fd_sc_hd__xnor2_1
X_5916_ _1836_ _1837_ _1839_ _1821_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__a31o_1
X_8635_ net221 _4082_ net220 vssd1 vssd1 vccd1 vccd1 _4086_ sky130_fd_sc_hd__a21oi_1
X_6896_ allocation.game.cactusDist.clock_div_inst0.counter\[0\] _2669_ _2671_ allocation.game.cactusDist.clock_div_inst0.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__or4b_1
XFILLER_0_14_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5847_ _1769_ _1770_ _1771_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__nand3_1
XFILLER_0_9_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5778_ _1699_ _1701_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8566_ net229 _3237_ vssd1 vssd1 vccd1 vccd1 _4017_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_12_clk_X clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4729_ _0645_ _0654_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__nand2_1
X_8497_ _3268_ _3282_ _3355_ _3271_ vssd1 vssd1 vccd1 vccd1 _3949_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_17_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7517_ allocation.game.lcdOutput.r_floor allocation.game.lcdOutput.r_cactus _3067_
+ _3070_ vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__nor4_1
XFILLER_0_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8684__A1 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7448_ _3059_ _3064_ _3018_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9042__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9090__RESET_B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7379_ _3010_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__inv_2
X_9118_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[12\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[12\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout87_A _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9049_ clknet_leaf_9_clk allocation.game.dinoJump.next_dinoY\[3\] net195 vssd1 vssd1
+ vccd1 vccd1 allocation.game.collision.dinoY\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__9192__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5670__A1 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8978__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5661__A1 _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7759__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6663__A _2516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6750_ allocation.game.cactus1size.clock_div_inst0.counter\[7\] _2573_ net158 vssd1
+ vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_34_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5701_ _1623_ _1625_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__nor2_1
XANTENNA__5964__A2 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6681_ allocation.game.lcdOutput.tft.spi.idle _0428_ net398 _2527_ vssd1 vssd1 vccd1
+ vccd1 _0104_ sky130_fd_sc_hd__a22o_1
XANTENNA__4911__A _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8902__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5632_ _1484_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__nor2_1
X_8420_ net115 _3871_ vssd1 vssd1 vccd1 vccd1 _3873_ sky130_fd_sc_hd__nor2_2
X_8351_ net140 _3809_ _3813_ vssd1 vssd1 vccd1 vccd1 _3814_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9065__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5563_ net72 _1435_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__nand2b_1
X_7302_ allocation.game.controller.init_module.delay_counter\[15\] allocation.game.controller.init_module.delay_counter\[14\]
+ allocation.game.controller.init_module.delay_counter\[13\] _2951_ vssd1 vssd1 vccd1
+ vccd1 _2957_ sky130_fd_sc_hd__and4_1
X_4514_ allocation.game.lcdOutput.framebufferIndex\[0\] net132 net130 vssd1 vssd1
+ vccd1 vccd1 _0453_ sky130_fd_sc_hd__and3_1
Xhold124 allocation.game.lcdOutput.tft.spi.internalSck vssd1 vssd1 vccd1 vccd1 net447
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 allocation.game.controller.init_module.delay_counter\[4\] vssd1 vssd1 vccd1
+ vccd1 net425 sky130_fd_sc_hd__dlygate4sd3_1
X_8282_ net81 _2260_ _2287_ net100 vssd1 vssd1 vccd1 vccd1 _3750_ sky130_fd_sc_hd__o22ai_1
Xhold113 allocation.game.cactus1size.clock_div_inst0.counter\[9\] vssd1 vssd1 vccd1
+ vccd1 net436 sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _1417_ _1418_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__and2_1
Xhold135 allocation.game.cactus2size.clock_div_inst1.counter\[6\] vssd1 vssd1 vccd1
+ vccd1 net458 sky130_fd_sc_hd__dlygate4sd3_1
X_7233_ allocation.game.dinoJump.count\[18\] _2905_ vssd1 vssd1 vccd1 vccd1 _2907_
+ sky130_fd_sc_hd__or2_1
Xhold146 allocation.game.controller.init_module.delay_counter\[1\] vssd1 vssd1 vccd1
+ vccd1 net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 allocation.game.cactusMove.x_dist\[1\] vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6397__X _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6838__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7164_ _2854_ _2853_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6115_ _2035_ _2038_ _2039_ _2012_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__a211oi_1
X_7095_ allocation.game.controller.drawBlock.x_start\[5\] _2772_ _2777_ allocation.game.controller.drawBlock.x_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__a22o_1
X_6046_ _1929_ _1944_ _1969_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__o21ai_1
X_7997_ _3490_ _3503_ _3505_ _3507_ vssd1 vssd1 vccd1 vccd1 _3508_ sky130_fd_sc_hd__a211o_1
X_6948_ _2399_ _2703_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__nor2_1
XANTENNA__4612__C1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9408__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6879_ net159 _2659_ _2660_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__nor3_1
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8618_ _4066_ _4067_ _4068_ vssd1 vssd1 vccd1 vccd1 _4069_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_49_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8549_ net217 net115 vssd1 vssd1 vccd1 vccd1 _4000_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6840__B1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9088__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5562__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7608__C1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7920_ allocation.game.controller.drawBlock.counter\[14\] allocation.game.controller.drawBlock.counter\[15\]
+ _3439_ allocation.game.controller.drawBlock.counter\[16\] vssd1 vssd1 vccd1 vccd1
+ _3446_ sky130_fd_sc_hd__a31o_1
X_7851_ net391 allocation.game.controller.drawBlock.state\[1\] allocation.game.controller.drawBlock.wr
+ _3399_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__a22o_1
X_6802_ allocation.game.cactus2size.clock_div_inst1.counter\[10\] _2606_ allocation.game.cactus2size.clock_div_inst1.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__a21oi_1
X_4994_ _0885_ _0887_ _0889_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__o21ai_1
X_7782_ net66 _3288_ net118 vssd1 vssd1 vccd1 vccd1 _3344_ sky130_fd_sc_hd__a21o_1
X_9521_ net306 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_6733_ allocation.game.cactus1size.clock_div_inst0.counter\[1\] allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6664_ _2517_ net228 _2515_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_pixel\[3\]
+ sky130_fd_sc_hd__mux2_1
X_9452_ clknet_leaf_18_clk _0359_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5737__A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9498__320 vssd1 vssd1 vccd1 vccd1 net320 _9498__320/LO sky130_fd_sc_hd__conb_1
X_8403_ net231 _3853_ vssd1 vssd1 vccd1 vccd1 _3858_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9029__RESET_B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5615_ _0769_ _0885_ _0887_ net88 vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9383_ clknet_leaf_13_clk net392 net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.wr
+ sky130_fd_sc_hd__dfstp_1
X_6595_ allocation.game.cactusMove.count\[7\] _2472_ _2474_ _2462_ vssd1 vssd1 vccd1
+ vccd1 allocation.game.cactusMove.n_count\[7\] sky130_fd_sc_hd__o211a_1
XFILLER_0_5_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8334_ net139 _3795_ _3796_ _3797_ vssd1 vssd1 vccd1 vccd1 _3798_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5546_ _1461_ _1463_ _1470_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__o21a_1
X_8265_ _2316_ _2317_ _2321_ vssd1 vssd1 vccd1 vccd1 _3736_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5477_ net64 _1355_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__or2_1
X_7216_ allocation.game.dinoJump.count\[12\] _2885_ _2893_ allocation.game.dinoJump.count\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__a31o_1
X_8196_ net282 _3684_ _3686_ vssd1 vssd1 vccd1 vccd1 _3687_ sky130_fd_sc_hd__or3b_1
X_7147_ _2848_ _2849_ _2847_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__a21o_1
X_7078_ allocation.game.controller.drawBlock.y_start\[2\] _2787_ _2795_ vssd1 vssd1
+ vccd1 vccd1 _2796_ sky130_fd_sc_hd__a21o_1
XANTENNA__6574__Y _2461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6029_ _1912_ _1952_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9230__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8327__B1 allocation.game.controller.drawBlock.y_end\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout63 _1053_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_4
Xfanout74 net76 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_4
Xfanout41 _3274_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout52 _3227_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_2
Xfanout85 _2863_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_1
XANTENNA__9380__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout96 net98 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_1_1__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6660__B _2461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7756__B net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload11 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinv_2
X_6380_ net280 allocation.game.cactusHeight1\[0\] _2290_ _2303_ vssd1 vssd1 vccd1
+ vccd1 _2304_ sky130_fd_sc_hd__a211oi_1
X_5400_ net61 _1324_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5331_ net65 _1255_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8050_ net265 net163 _3556_ _3558_ _3553_ vssd1 vssd1 vccd1 vccd1 _3559_ sky130_fd_sc_hd__a221o_1
XANTENNA__9103__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5855__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5262_ _1183_ _1185_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__or2_1
X_7001_ _2736_ _2737_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__nor2_1
X_5193_ _1114_ _1116_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9253__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8952_ net116 _3704_ vssd1 vssd1 vccd1 vccd1 _4401_ sky130_fd_sc_hd__nand2_1
X_7903_ allocation.game.controller.drawBlock.counter\[10\] allocation.game.controller.drawBlock.counter\[11\]
+ _3430_ vssd1 vssd1 vccd1 vccd1 _3434_ sky130_fd_sc_hd__and3_1
X_8883_ _3866_ _3874_ _3876_ vssd1 vssd1 vccd1 vccd1 _4333_ sky130_fd_sc_hd__o21a_1
X_7834_ _3391_ _3384_ _2367_ vssd1 vssd1 vccd1 vccd1 _3392_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7765_ _3299_ _3324_ vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4977_ _0594_ _0698_ _0699_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__a21oi_2
XANTENNA__5467__A _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6716_ allocation.game.cactus1size.clock_div_inst1.counter\[10\] _2549_ _2551_ vssd1
+ vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__o21a_1
X_9504_ net289 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4802__C _0708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload5/X sky130_fd_sc_hd__clkbuf_4
X_7696_ _3252_ _3257_ vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__nor2_1
X_9435_ clknet_leaf_11_clk _0344_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6647_ allocation.game.cactusMove.count\[27\] _2506_ vssd1 vssd1 vccd1 vccd1 _2507_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6578_ net147 _2452_ _2463_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[1\]
+ sky130_fd_sc_hd__and3_1
X_9366_ clknet_leaf_4_clk _0015_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.bcd_tens\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8317_ net275 _3472_ _3522_ vssd1 vssd1 vccd1 vccd1 _3782_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5529_ _1453_ _1452_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__and2b_1
X_9297_ clknet_leaf_21_clk _0083_ net180 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5846__A1 _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8248_ _3000_ _3724_ _3035_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__o21ai_1
Xfanout231 allocation.game.controller.v\[6\] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_4
Xfanout220 allocation.game.cactusMove.pixel\[7\] vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
X_8179_ _0642_ _0643_ _0656_ vssd1 vssd1 vccd1 vccd1 _3671_ sky130_fd_sc_hd__and3_1
XANTENNA__5846__B2 _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 allocation.game.controller.state\[8\] vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
Xfanout264 net267 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout253 allocation.game.lcdOutput.tft.initSeqCounter\[0\] vssd1 vssd1 vccd1 vccd1
+ net253 sky130_fd_sc_hd__buf_2
XANTENNA__4817__Y _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 allocation.game.collision.dinoY\[2\] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7220__B1 _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9126__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9276__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8787__B1 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4900_ _0823_ _0824_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5880_ _1764_ _1802_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4831_ _0737_ _0755_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4762_ _0642_ _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__and2b_1
X_7550_ _3152_ _3153_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__and2_1
X_6501_ _2409_ _2410_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__or2_1
X_4693_ net226 net224 _0619_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7481_ _3047_ _3052_ net249 vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6432_ _2354_ allocation.game.game.score\[2\] _2320_ vssd1 vssd1 vccd1 vccd1 _2355_
+ sky130_fd_sc_hd__mux2_1
X_9220_ clknet_leaf_22_clk _0046_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_9151_ clknet_leaf_20_clk _0215_ net199 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.x_dist\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6363_ _2278_ _2286_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__nand2_1
X_8102_ _0654_ _0682_ _2406_ _3603_ vssd1 vssd1 vccd1 vccd1 _3605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9082_ clknet_leaf_14_clk _0178_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_5314_ _1238_ _1236_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__and2b_1
X_6294_ _0432_ _2185_ _2187_ allocation.game.controller.drawBlock.counter\[10\] _2218_
+ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__o221a_1
X_5245_ _1052_ _1113_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__xnor2_1
X_8033_ _3541_ vssd1 vssd1 vccd1 vccd1 _3542_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold28 _0248_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 allocation.game.lcdOutput.tft.spi.dataShift\[3\] vssd1 vssd1 vccd1 vccd1 net340
+ sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _1099_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__or2_1
Xhold39 _0255_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8935_ _0462_ net199 _4384_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8866_ _4454_ net275 vssd1 vssd1 vccd1 vccd1 _4316_ sky130_fd_sc_hd__and2_1
X_7817_ _2353_ _3376_ vssd1 vssd1 vccd1 vccd1 _3377_ sky130_fd_sc_hd__xnor2_1
X_8797_ _4231_ _4233_ vssd1 vssd1 vccd1 vccd1 _4247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9149__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7748_ _3304_ _3309_ _3307_ vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__a21bo_1
X_7679_ _3230_ _3235_ _3232_ vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__a21oi_1
X_9418_ clknet_leaf_13_clk _0327_ net210 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.idx\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8702__B1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9299__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9349_ clknet_leaf_1_clk _0281_ net165 vssd1 vssd1 vccd1 vccd1 allocation.game.bcd_ones\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__8955__B _3256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6492__A1 _0417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout72_X net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8211__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5030_ _0946_ _0953_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__xor2_1
XANTENNA__6666__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6981_ _2724_ net92 _2723_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__and3b_1
X_5932_ _1854_ _1855_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__xnor2_1
X_8720_ net257 _3249_ _4141_ _4166_ vssd1 vssd1 vccd1 vccd1 _4171_ sky130_fd_sc_hd__a31o_1
XANTENNA__4633__B allocation.game.controller.drawBlock.x_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_5863_ _1784_ _1787_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__nand2_1
X_8651_ net111 net76 vssd1 vssd1 vccd1 vccd1 _4102_ sky130_fd_sc_hd__nor2_1
X_4814_ _0710_ net103 vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__or2_2
X_8582_ _0613_ _2375_ net219 vssd1 vssd1 vccd1 vccd1 _4033_ sky130_fd_sc_hd__a21o_1
X_5794_ _1671_ _1673_ _1672_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__a21o_1
X_7602_ allocation.game.cactusDist.clock_div_inst1.clk1 allocation.game.cactusDist.lfsr2\[0\]
+ allocation.game.cactusDist.lfsr2\[1\] net143 vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__a31o_1
X_4745_ _0665_ _0667_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__xnor2_2
X_7533_ _3078_ _3083_ net249 vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5745__A _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4676_ net236 _0575_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7464_ net250 _3076_ _3079_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__o21ai_1
X_7395_ allocation.game.controller.color\[11\] net203 _3016_ _3017_ vssd1 vssd1 vccd1
+ vccd1 _0219_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6415_ _2328_ _2335_ _2337_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9203_ _0141_ _0413_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6346_ allocation.game.collision.dinoY\[0\] allocation.game.cactusHeight2\[0\] vssd1
+ vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__nand2_1
X_9134_ clknet_leaf_2_clk allocation.game.cactusMove.n_count\[28\] net176 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[28\] sky130_fd_sc_hd__dfrtp_1
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
X_9065_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[11\] net192 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8016_ net135 _3520_ _3524_ _3525_ vssd1 vssd1 vccd1 vccd1 _3526_ sky130_fd_sc_hd__a31o_1
X_6277_ _2095_ _2201_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__nand2_1
X_5228_ _1143_ _1146_ net60 vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__a21o_1
X_5159_ _1082_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8918_ net38 _4367_ vssd1 vssd1 vccd1 vccd1 _4368_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8849_ allocation.game.lcdOutput.framebufferIndex\[0\] net280 vssd1 vssd1 vccd1 vccd1
+ _4299_ sky130_fd_sc_hd__xor2_1
XANTENNA__7694__X _3256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8975__A2_N net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9314__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9464__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4530_ net264 net261 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7180_ _0471_ _2867_ _2869_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6200_ _1424_ _2123_ _1422_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__a21o_1
X_6131_ net110 _0900_ _2055_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6062_ _0723_ _0904_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__nor2_1
X_5013_ _0772_ _0831_ _0866_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__a21o_1
XANTENNA__7956__A1 allocation.game.controller.drawBlock.y_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6964_ allocation.game.scoreCounter.clock_div.counter\[12\] _2712_ net93 vssd1 vssd1
+ vccd1 vccd1 _2714_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_18_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6895_ allocation.game.cactusDist.clock_div_inst0.counter\[11\] allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ allocation.game.cactusDist.clock_div_inst0.counter\[13\] allocation.game.cactusDist.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__or4_1
X_5915_ _1836_ _1837_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__nand3_1
X_8703_ _4152_ _4153_ vssd1 vssd1 vccd1 vccd1 _4154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8634_ _3997_ _4000_ _4084_ vssd1 vssd1 vccd1 vccd1 _4085_ sky130_fd_sc_hd__a21oi_1
X_5846_ _0722_ _0885_ _0887_ _0716_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8565_ _4013_ _4014_ _4015_ vssd1 vssd1 vccd1 vccd1 _4016_ sky130_fd_sc_hd__and3_1
X_5777_ _1699_ _1701_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7516_ _3020_ _3127_ vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8496_ net56 _3298_ _3328_ _3871_ vssd1 vssd1 vccd1 vccd1 _3948_ sky130_fd_sc_hd__and4_1
X_4728_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4659_ _0587_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__nand2b_1
X_7447_ _3044_ _3049_ _3050_ _3063_ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__a31o_1
X_7378_ _3009_ _3008_ vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_10_Left_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9117_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[11\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[11\] sky130_fd_sc_hd__dfrtp_1
X_6329_ allocation.game.cactusHeight2\[3\] _2238_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__xnor2_2
XANTENNA__9337__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6447__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9048_ clknet_leaf_3_clk allocation.game.dinoJump.next_dinoY\[2\] net193 vssd1 vssd1
+ vccd1 vccd1 allocation.game.collision.dinoY\[2\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9406__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9487__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5700_ _0762_ _0886_ _0888_ _0738_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__o22a_1
XANTENNA__7775__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6680_ allocation.game.lcdOutput.tft.spi.counter\[2\] allocation.game.lcdOutput.tft.spi.counter\[1\]
+ _2526_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__and3_1
XANTENNA__4470__Y _4459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5631_ _0732_ _1483_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__nor2_1
X_8350_ net136 _3810_ _3812_ _3556_ vssd1 vssd1 vccd1 vccd1 _3813_ sky130_fd_sc_hd__o31a_1
X_5562_ net82 _1486_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__nand2_1
X_7301_ allocation.game.controller.init_module.delay_counter\[14\] _2951_ _2955_ vssd1
+ vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8281_ net244 _3746_ _3748_ _3481_ vssd1 vssd1 vccd1 vccd1 _3749_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4513_ allocation.game.lcdOutput.framebufferIndex\[0\] net132 net130 vssd1 vssd1
+ vccd1 vccd1 _0452_ sky130_fd_sc_hd__a21oi_1
Xhold125 allocation.game.dinoJump.count\[14\] vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__dlygate4sd3_1
X_7232_ net84 _2904_ _2906_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__and3_1
Xhold103 allocation.game.cactusHeight2\[2\] vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 allocation.game.cactusDist.clock_div_inst1.counter\[12\] vssd1 vssd1 vccd1
+ vccd1 net437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5493_ _1411_ _1415_ _1416_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__or3_1
Xhold158 allocation.game.cactusMove.count\[4\] vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold147 allocation.game.controller.init_module.delay_counter\[3\] vssd1 vssd1 vccd1
+ vccd1 net470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold136 allocation.game.cactus2size.clock_div_inst0.counter\[12\] vssd1 vssd1 vccd1
+ vccd1 net459 sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ _2850_ _2852_ _2855_ _2845_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7094_ allocation.game.controller.color\[10\] _2792_ _2803_ vssd1 vssd1 vccd1 vccd1
+ _2809_ sky130_fd_sc_hd__a21o_1
X_6114_ _2009_ _2011_ _2010_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__a21oi_1
X_6045_ _1929_ _1944_ _1969_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7996_ _3506_ vssd1 vssd1 vccd1 vccd1 _3507_ sky130_fd_sc_hd__inv_2
X_6947_ allocation.game.scoreCounter.clock_div.counter\[6\] _2398_ net91 vssd1 vssd1
+ vccd1 vccd1 _2703_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6878_ allocation.game.cactusDist.clock_div_inst1.counter\[7\] allocation.game.cactusDist.clock_div_inst1.counter\[8\]
+ _2656_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5829_ _1752_ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8617_ net97 _4065_ vssd1 vssd1 vccd1 vccd1 _4068_ sky130_fd_sc_hd__or2_1
X_8548_ net217 net115 vssd1 vssd1 vccd1 vccd1 _3999_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5933__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8479_ _3915_ _3931_ vssd1 vssd1 vccd1 vccd1 _3932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4836__X _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8593__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4603__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5843__A _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9328__RESET_B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_11_clk_X clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7850_ net236 allocation.game.controller.drawBlock.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _3399_ sky130_fd_sc_hd__nand2_1
XANTENNA__7387__A2 _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6801_ allocation.game.cactus2size.clock_div_inst1.counter\[10\] _2606_ _2608_ vssd1
+ vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__o21a_1
XANTENNA__9032__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4993_ net79 net86 vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__nor2_1
X_7781_ net34 net40 _3313_ _3342_ vssd1 vssd1 vccd1 vccd1 _3343_ sky130_fd_sc_hd__o22a_1
X_9520_ net305 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
X_6732_ allocation.game.cactus1size.clock_div_inst0.counter\[1\] allocation.game.cactus1size.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6663_ _2516_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9451_ clknet_leaf_18_clk _0358_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8402_ net231 _3853_ vssd1 vssd1 vccd1 vccd1 _3857_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5614_ _0777_ _0892_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6594_ allocation.game.cactusMove.count\[7\] _2472_ vssd1 vssd1 vccd1 vccd1 _2474_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9382_ clknet_leaf_3_clk _0292_ net199 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight2\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8333_ net139 _3794_ _3556_ vssd1 vssd1 vccd1 vccd1 _3797_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5545_ _1468_ _1469_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__nor2_1
X_8264_ allocation.game.game.score\[2\] allocation.game.game.score\[1\] allocation.game.game.score\[4\]
+ allocation.game.game.score\[3\] vssd1 vssd1 vccd1 vccd1 _3735_ sky130_fd_sc_hd__a211oi_1
X_5476_ net64 _1400_ _1399_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__a21o_1
X_7215_ allocation.game.dinoJump.count\[12\] _2891_ _2894_ net84 vssd1 vssd1 vccd1
+ vccd1 _0162_ sky130_fd_sc_hd__o211a_1
X_8195_ _2373_ _2375_ net100 _3685_ vssd1 vssd1 vccd1 vccd1 _3686_ sky130_fd_sc_hd__a211o_1
X_7146_ allocation.game.lcdOutput.framebufferIndex\[11\] _2838_ vssd1 vssd1 vccd1
+ vccd1 _2849_ sky130_fd_sc_hd__nand2_1
XANTENNA_input4_A gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7077_ allocation.game.controller.drawBlock.x_start\[2\] _2772_ _2777_ allocation.game.controller.drawBlock.x_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__a22o_1
X_6028_ _1909_ _1911_ _1910_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__a21o_1
XANTENNA__7686__Y _3248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7979_ net137 _3489_ _3490_ _3487_ _3488_ vssd1 vssd1 vccd1 vccd1 _3491_ sky130_fd_sc_hd__a32o_1
XANTENNA__8304__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout53 _0233_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_2
Xfanout42 _3267_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_2
Xfanout64 net65 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_4
Xfanout97 net98 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout86 _0891_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_4
Xfanout75 net76 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9055__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5557__B _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload12 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload12/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__6669__A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _1253_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__and2_1
X_5261_ _1183_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7000_ allocation.game.bcd_ones\[1\] allocation.game.bcd_ones\[2\] vssd1 vssd1 vccd1
+ vccd1 _2737_ sky130_fd_sc_hd__and2b_1
X_5192_ _1114_ _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4917__A _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8951_ net116 _3704_ vssd1 vssd1 vccd1 vccd1 _4400_ sky130_fd_sc_hd__or2_1
X_7902_ net94 _3432_ _3433_ net109 allocation.game.controller.drawBlock.counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__a32o_1
X_8882_ _3299_ _3919_ vssd1 vssd1 vccd1 vccd1 _4332_ sky130_fd_sc_hd__nor2_1
X_7833_ _2361_ _2367_ _3390_ _2348_ _2343_ vssd1 vssd1 vccd1 vccd1 _3391_ sky130_fd_sc_hd__o32a_1
XFILLER_0_4_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7764_ _3324_ _3325_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4976_ net78 net124 vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__nor2_2
X_6715_ allocation.game.cactus1size.clock_div_inst1.counter\[10\] _2549_ net158 vssd1
+ vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__a21oi_1
X_9503_ net288 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
X_7695_ allocation.game.lcdOutput.framebufferIndex\[4\] net46 vssd1 vssd1 vccd1 vccd1
+ _3257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload6 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload6/X sky130_fd_sc_hd__clkbuf_4
X_9434_ clknet_leaf_11_clk _0343_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_6646_ _2506_ net150 _2505_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[26\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8778__B _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6577_ allocation.game.cactusMove.count\[1\] allocation.game.cactusMove.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__nand2_1
X_9365_ clknet_leaf_5_clk _0014_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.bcd_tens\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_8316_ _3529_ _3767_ _3779_ _3780_ net135 vssd1 vssd1 vccd1 vccd1 _3781_ sky130_fd_sc_hd__o311a_1
XFILLER_0_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5528_ _0792_ _1440_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__xnor2_1
X_9296_ clknet_leaf_21_clk _0082_ net180 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5459_ _1333_ _1383_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__and2_1
XANTENNA__8794__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8247_ allocation.game.lcdOutput.tft.remainingDelayTicks\[13\] _2991_ vssd1 vssd1
+ vccd1 vccd1 _3724_ sky130_fd_sc_hd__xor2_1
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
XANTENNA__9078__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout221 net223 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
X_8178_ net121 _3667_ vssd1 vssd1 vccd1 vccd1 _3670_ sky130_fd_sc_hd__and2b_1
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5846__A2 _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout243 allocation.game.controller.state\[1\] vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
Xfanout265 net267 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
X_7129_ allocation.game.lcdOutput.framebufferIndex\[7\] allocation.game.lcdOutput.framebufferIndex\[8\]
+ _2832_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__and3_1
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_4
Xfanout276 allocation.game.collision.dinoY\[2\] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8796__A1 _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout62_A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8034__A allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5658__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8720__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5534__A1 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4737__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4830_ _0552_ _0569_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_16_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4761_ net142 _0686_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6500_ allocation.game.controller.state\[6\] net243 net238 vssd1 vssd1 vccd1 vccd1
+ _2410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4692_ net226 _0619_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7480_ _3042_ _3074_ _3093_ net248 vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6431_ _2322_ _2329_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__or2_1
X_6362_ allocation.game.cactusHeight1\[1\] allocation.game.cactusHeight1\[0\] vssd1
+ vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__or2_1
X_9150_ clknet_leaf_3_clk _0214_ net199 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.x_dist\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8101_ net228 net101 _2516_ allocation.game.controller.state\[2\] vssd1 vssd1 vccd1
+ vccd1 _3604_ sky130_fd_sc_hd__a2bb2o_1
X_5313_ _1030_ _1237_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__xnor2_1
X_9081_ clknet_leaf_14_clk _0177_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6293_ allocation.game.controller.drawBlock.counter\[10\] _2187_ _2188_ allocation.game.controller.drawBlock.counter\[9\]
+ _2217_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__a221oi_1
XANTENNA__9220__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5244_ net62 _1168_ _1166_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__a21o_1
X_8032_ _3539_ _3540_ vssd1 vssd1 vccd1 vccd1 _3541_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5175_ _0924_ _1098_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__and2_1
Xhold18 _0245_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 allocation.game.cactus2size.clock_div_inst1.counter\[13\] vssd1 vssd1 vccd1
+ vccd1 net352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9370__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8934_ _4276_ _4302_ _4334_ _4294_ _4383_ vssd1 vssd1 vccd1 vccd1 _4384_ sky130_fd_sc_hd__a221o_1
XANTENNA__6581__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8865_ net272 net128 vssd1 vssd1 vccd1 vccd1 _4315_ sky130_fd_sc_hd__or2_1
XANTENNA__7677__B net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7816_ _2360_ _2385_ _2370_ vssd1 vssd1 vccd1 vccd1 _3376_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_17_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8950__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8796_ _3770_ _4225_ _0442_ vssd1 vssd1 vccd1 vccd1 _4246_ sky130_fd_sc_hd__a21oi_1
X_4959_ _0854_ _0883_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7747_ _3308_ net50 _3237_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__and3b_1
XFILLER_0_35_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7678_ allocation.game.lcdOutput.framebufferIndex\[6\] _3229_ net48 vssd1 vssd1 vccd1
+ vccd1 _3240_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9417_ clknet_leaf_13_clk _0326_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.idx\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6629_ allocation.game.cactusMove.count\[19\] allocation.game.cactusMove.count\[20\]
+ _2492_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__and3_1
XANTENNA__8702__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9348_ clknet_leaf_20_clk _0280_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.r_win
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9279_ clknet_leaf_1_clk _0090_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5941__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout65_X net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4844__X _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7868__A allocation.game.controller.drawBlock.state\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8699__A _3208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9243__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9393__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5570__B _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6980_ allocation.game.scoreCounter.clock_div.counter\[18\] allocation.game.scoreCounter.clock_div.counter\[17\]
+ _2721_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__and3_1
X_5931_ _1854_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5862_ _1784_ _1785_ _1786_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8650_ net111 net76 vssd1 vssd1 vccd1 vccd1 _4101_ sky130_fd_sc_hd__nand2_1
X_4813_ _0735_ _0736_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8581_ _3997_ _4031_ _3999_ vssd1 vssd1 vccd1 vccd1 _4032_ sky130_fd_sc_hd__a21o_1
X_7601_ allocation.game.cactusDist.clock_div_inst1.clk1 allocation.game.cactusDist.lfsr2\[1\]
+ allocation.game.cactusDist.lfsr2\[0\] vssd1 vssd1 vccd1 vccd1 _3173_ sky130_fd_sc_hd__a21oi_1
X_5793_ _1714_ _1716_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__xor2_1
XANTENNA__8402__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4930__A _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7532_ net367 net53 _3129_ _3141_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4744_ _0669_ _0670_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5745__B _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4675_ _0602_ _0603_ _0576_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__a21o_2
XFILLER_0_25_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9202_ _0140_ _0412_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_7463_ _3058_ _3078_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__and2_1
X_7394_ net239 _2381_ _2409_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__a21o_1
X_6414_ allocation.game.game.score\[5\] _2324_ _2336_ vssd1 vssd1 vccd1 vccd1 _2337_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6345_ _2244_ _2266_ _2267_ _2268_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__and4_1
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
X_9133_ clknet_leaf_2_clk allocation.game.cactusMove.n_count\[27\] net176 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9064_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[10\] net192 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6276_ _2092_ _2094_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__or2_1
X_5227_ _1150_ _1151_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__or2_1
X_8015_ _0504_ _3518_ _3519_ net138 vssd1 vssd1 vccd1 vccd1 _3525_ sky130_fd_sc_hd__o211a_1
X_5158_ _1077_ _1079_ _1081_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__or3b_1
X_5089_ _1002_ _1003_ _0999_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__a21o_1
XANTENNA__9116__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8917_ net258 _4364_ vssd1 vssd1 vccd1 vccd1 _4367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8848_ _4297_ vssd1 vssd1 vccd1 vccd1 _4298_ sky130_fd_sc_hd__inv_2
XANTENNA__9265__RESET_B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9266__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8779_ _4226_ _4228_ vssd1 vssd1 vccd1 vccd1 _4229_ sky130_fd_sc_hd__or2_1
XANTENNA__8031__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6465__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7780__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6130_ _1946_ _2019_ _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6061_ net141 net102 _1947_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__or3_1
X_5012_ _0935_ _0936_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6963_ allocation.game.scoreCounter.clock_div.counter\[12\] _2712_ vssd1 vssd1 vccd1
+ vccd1 _2713_ sky130_fd_sc_hd__and2_1
XANTENNA__9289__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6894_ allocation.game.cactusDist.clock_div_inst0.counter\[7\] allocation.game.cactusDist.clock_div_inst0.counter\[6\]
+ allocation.game.cactusDist.clock_div_inst0.counter\[9\] allocation.game.cactusDist.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8702_ net104 _4151_ net89 vssd1 vssd1 vccd1 vccd1 _4153_ sky130_fd_sc_hd__a21o_1
X_5914_ _1776_ _1838_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8633_ net221 net220 _4082_ vssd1 vssd1 vccd1 vccd1 _4084_ sky130_fd_sc_hd__and3_1
X_5845_ _0741_ net86 vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5195__A2 _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8564_ net68 _3676_ vssd1 vssd1 vccd1 vccd1 _4015_ sky130_fd_sc_hd__or2_1
X_5776_ _1648_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__and2_1
X_4727_ _0636_ _0653_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__or2_2
X_8495_ _3295_ _3297_ _3880_ vssd1 vssd1 vccd1 vccd1 _3947_ sky130_fd_sc_hd__o21ai_1
X_7515_ _3021_ _3077_ _3124_ _3126_ vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__o211a_1
X_4658_ allocation.game.controller.drawBlock.y_end\[2\] allocation.game.controller.drawBlock.y_start\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7446_ _3051_ _3060_ _3061_ _3062_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8278__S net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7690__B net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4589_ _4456_ allocation.game.controller.v\[0\] vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__nand2_2
X_9116_ clknet_leaf_6_clk allocation.game.cactusMove.n_count\[10\] net172 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[10\] sky130_fd_sc_hd__dfrtp_1
X_7377_ allocation.game.cactusDist.lfsr1\[0\] allocation.game.cactusDist.lfsr2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__xnor2_2
X_6328_ net271 _2249_ _2251_ _2247_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__o211a_1
XANTENNA__4819__B _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9047_ clknet_leaf_9_clk allocation.game.dinoJump.next_dinoY\[1\] net195 vssd1 vssd1
+ vccd1 vccd1 allocation.game.collision.dinoY\[1\] sky130_fd_sc_hd__dfrtp_1
X_6259_ allocation.game.controller.drawBlock.counter\[12\] _2183_ vssd1 vssd1 vccd1
+ vccd1 _2184_ sky130_fd_sc_hd__nand2_1
XANTENNA__9446__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4570__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8109__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9431__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8060__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7775__B net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7571__B1 _2526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6374__A1 _4459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5630_ net72 _1554_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__and2_1
X_5561_ _1481_ _1484_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__xnor2_1
X_7300_ allocation.game.controller.init_module.delay_counter\[14\] allocation.game.controller.init_module.delay_counter\[13\]
+ _2951_ vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__and3_1
X_8280_ net137 _3482_ _3747_ _3473_ net241 vssd1 vssd1 vccd1 vccd1 _3748_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4512_ net255 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__inv_2
X_5492_ _1411_ _1415_ _1416_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__o21ai_1
Xhold104 allocation.game.controller.drawBlock.y_start\[3\] vssd1 vssd1 vccd1 vccd1
+ net427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6678__Y _2526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7231_ _2905_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__inv_2
Xhold126 allocation.game.controller.drawBlock.x_start\[8\] vssd1 vssd1 vccd1 vccd1
+ net449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold115 allocation.game.cactus2size.clock_div_inst1.clk1 vssd1 vssd1 vccd1 vccd1
+ net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 allocation.game.controller.init_module.delay_counter\[16\] vssd1 vssd1 vccd1
+ vccd1 net460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold148 allocation.game.dinoJump.dinoDelay\[19\] vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 allocation.game.cactus2size.clock_div_inst0.counter\[6\] vssd1 vssd1 vccd1
+ vccd1 net482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7162_ _2852_ _2860_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__xor2_1
X_7093_ _2759_ _2789_ _2807_ _2808_ vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__o22a_1
XANTENNA_clkload14_A clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6113_ _2035_ _2036_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__nand3_1
X_6044_ net141 _0730_ _1967_ _1968_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7995_ _0490_ _3490_ vssd1 vssd1 vccd1 vccd1 _3506_ sky130_fd_sc_hd__or2_1
X_6946_ _2398_ net91 _2702_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9046__SET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6877_ allocation.game.cactusDist.clock_div_inst1.counter\[7\] _2656_ allocation.game.cactusDist.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5828_ _0732_ _1120_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__xnor2_1
X_8616_ net119 _4063_ vssd1 vssd1 vccd1 vccd1 _4067_ sky130_fd_sc_hd__or2_1
X_5759_ _0770_ _0778_ _0906_ _0908_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__or4_1
X_8547_ _3997_ vssd1 vssd1 vccd1 vccd1 _3998_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5933__B net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9304__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8478_ net119 net50 _3866_ _3882_ _3876_ vssd1 vssd1 vccd1 vccd1 _3931_ sky130_fd_sc_hd__a41o_1
X_7429_ allocation.game.lcdOutput.tft.initSeqCounter\[0\] net252 vssd1 vssd1 vccd1
+ vccd1 _3046_ sky130_fd_sc_hd__and2_1
XANTENNA__5013__X _0938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5843__B _0886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6020__A _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8281__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4746__Y _0673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6800_ allocation.game.cactus2size.clock_div_inst1.counter\[10\] _2606_ net162 vssd1
+ vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7780_ _2827_ net34 _3341_ vssd1 vssd1 vccd1 vccd1 _3342_ sky130_fd_sc_hd__or3b_1
X_4992_ _0897_ _0916_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__xnor2_2
X_6731_ allocation.game.cactus1size.clock_div_inst0.counter\[0\] net154 _2561_ vssd1
+ vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__and3b_1
XANTENNA__9327__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9450_ clknet_leaf_18_clk _0357_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6662_ _0611_ _0619_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__or2_2
X_8401_ net231 net85 vssd1 vssd1 vccd1 vccd1 _3856_ sky130_fd_sc_hd__nand2_1
X_5613_ net87 _0885_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__and2_1
X_9381_ clknet_leaf_10_clk _0291_ net196 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8332_ net265 _3782_ vssd1 vssd1 vccd1 vccd1 _3796_ sky130_fd_sc_hd__nand2_1
X_6593_ _2472_ _2473_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5544_ _1409_ _1467_ _1465_ _1437_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_48_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9477__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8263_ _3034_ _3734_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__or2_1
X_5475_ _1397_ _1398_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__xnor2_1
X_7214_ allocation.game.dinoJump.count\[12\] _2891_ vssd1 vssd1 vccd1 vccd1 _2894_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8194_ allocation.game.cactusMove.pixel\[5\] _2373_ net223 vssd1 vssd1 vccd1 vccd1
+ _3685_ sky130_fd_sc_hd__a21oi_1
X_7145_ allocation.game.lcdOutput.framebufferIndex\[12\] _2839_ vssd1 vssd1 vccd1
+ vccd1 _2848_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7076_ _2791_ _2793_ _2794_ _2789_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__o31a_1
X_6027_ _1949_ _1950_ _1948_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_1_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7978_ _0494_ _3470_ _0500_ vssd1 vssd1 vccd1 vccd1 _3490_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_25_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ allocation.game.cactusDist.clock_div_inst0.counter\[11\] allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ _2690_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout54 net55 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout65 _0917_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_4
Xfanout43 _3267_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_2
Xfanout87 _0759_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_2
Xfanout76 _3199_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_4
Xfanout98 _3191_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5854__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload13 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_4
XANTENNA__6669__B _2461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5260_ _1140_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5191_ _1055_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8950_ net69 _3673_ _4396_ _4398_ vssd1 vssd1 vccd1 vccd1 _4399_ sky130_fd_sc_hd__a211o_1
XANTENNA__8006__A1 _3516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7901_ allocation.game.controller.drawBlock.counter\[10\] _3430_ vssd1 vssd1 vccd1
+ vccd1 _3433_ sky130_fd_sc_hd__or2_1
X_8881_ net258 _0467_ _4326_ _4330_ vssd1 vssd1 vccd1 vccd1 _4331_ sky130_fd_sc_hd__a22o_1
XANTENNA__4933__A _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7832_ _3388_ _3389_ _3387_ vssd1 vssd1 vccd1 vccd1 _3390_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9380__SET_B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4975_ net124 vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__inv_2
X_7763_ net114 _3302_ vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6714_ _2549_ _2550_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__nor2_1
X_9502_ net287 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
X_9433_ clknet_leaf_11_clk _0342_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_7694_ _3254_ _3255_ vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload7 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__clkinv_8
X_6645_ allocation.game.cactusMove.count\[25\] allocation.game.cactusMove.count\[26\]
+ _2502_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6576_ allocation.game.cactusMove.count\[0\] _2462_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[0\]
+ sky130_fd_sc_hd__and2b_1
XANTENNA__8140__A _0673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9364_ clknet_leaf_4_clk _0013_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.bcd_tens\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8315_ _3529_ _3767_ _3779_ vssd1 vssd1 vccd1 vccd1 _3780_ sky130_fd_sc_hd__o21ai_1
X_5527_ _0838_ _1196_ _1443_ _1451_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__a31o_1
X_9295_ clknet_leaf_21_clk _0081_ net189 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_8246_ _3027_ _3723_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__nand2_1
X_5458_ _1331_ _1332_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout200 allocation.game.cactus1size.clock_div_inst0.reset vssd1 vssd1 vccd1 vccd1
+ net200 sky130_fd_sc_hd__clkbuf_4
Xfanout211 net215 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_2
X_8177_ _3666_ _3669_ allocation.game.controller.drawBlock.x_start\[4\] net205 vssd1
+ vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__o2bb2a_1
X_5389_ _1296_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout244 allocation.game.controller.state\[4\] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
Xfanout233 allocation.game.cactus1size.state\[1\] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_4
X_7128_ allocation.game.lcdOutput.framebufferIndex\[7\] _2832_ vssd1 vssd1 vccd1 vccd1
+ _0412_ sky130_fd_sc_hd__xor2_1
Xfanout255 allocation.game.lcdOutput.tft.frameBufferLowNibble vssd1 vssd1 vccd1 vccd1
+ net255 sky130_fd_sc_hd__clkbuf_8
X_7059_ _2774_ _2778_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__nor2_2
Xfanout277 allocation.game.collision.dinoY\[2\] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_2
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5939__A _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5658__B _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4990__B1 net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_clk_X clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6495__B1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4760_ net142 _0655_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4691_ net230 net227 vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7783__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6430_ _2328_ _2351_ _2352_ _2319_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_45_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6361_ net273 _2280_ _2281_ _2283_ _2284_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5312_ _1179_ _1180_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__xor2_1
X_8100_ _0686_ _3602_ vssd1 vssd1 vccd1 vccd1 _3603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8895__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9080_ clknet_leaf_14_clk _0176_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6292_ allocation.game.controller.drawBlock.counter\[9\] _2188_ _2216_ vssd1 vssd1
+ vccd1 vccd1 _2217_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5243_ _1166_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__nor2_1
X_8031_ allocation.game.collision.dinoY\[3\] net270 net266 vssd1 vssd1 vccd1 vccd1
+ _3540_ sky130_fd_sc_hd__and3_2
X_5174_ _0924_ _1098_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__nor2_1
Xhold19 allocation.game.cactusDist.clock_div_inst0.counter\[13\] vssd1 vssd1 vccd1
+ vccd1 net342 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4647__B allocation.game.controller.drawBlock.y_end\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8933_ _4215_ _4336_ _4339_ _4341_ _4382_ vssd1 vssd1 vccd1 vccd1 _4383_ sky130_fd_sc_hd__a41o_1
X_8864_ net272 net128 vssd1 vssd1 vccd1 vccd1 _4314_ sky130_fd_sc_hd__nand2_1
X_7815_ _3177_ _3375_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__nand2_1
XANTENNA__7974__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8795_ _0468_ _4243_ vssd1 vssd1 vccd1 vccd1 _4245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4958_ _0863_ _0881_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7746_ _3249_ net46 vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__or2_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4889_ _0806_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7677_ allocation.game.lcdOutput.framebufferIndex\[6\] net48 vssd1 vssd1 vccd1 vccd1
+ _3239_ sky130_fd_sc_hd__xor2_4
X_9416_ clknet_leaf_13_clk _0325_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.idx\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6628_ allocation.game.cactusMove.count\[19\] allocation.game.cactusMove.count\[18\]
+ _2490_ allocation.game.cactusMove.count\[20\] vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9045__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9347_ clknet_leaf_4_clk _0279_ net173 vssd1 vssd1 vccd1 vccd1 allocation.game.game.score\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_6559_ allocation.game.dinoJump.dinoDelay\[19\] _2447_ vssd1 vssd1 vccd1 vccd1 _2448_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9278_ clknet_leaf_3_clk _0266_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.clk1
+ sky130_fd_sc_hd__dfxtp_1
X_8229_ _2987_ _3712_ vssd1 vssd1 vccd1 vccd1 _3713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4748__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7968__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6640__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5930_ _1804_ _1805_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__xnor2_1
X_5861_ _1735_ _1783_ _1782_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__a21o_1
X_7600_ net143 _3172_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__or2_1
X_4812_ _0735_ _0736_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__and2_4
X_8580_ _0613_ _2524_ vssd1 vssd1 vccd1 vccd1 _4031_ sky130_fd_sc_hd__nand2_1
X_5792_ _1716_ _1714_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7531_ _0233_ _3140_ vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__nand2_1
XANTENNA__9068__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4743_ net217 _0664_ _0668_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7462_ net252 _3054_ vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__or2_1
X_4674_ _0576_ _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6413_ allocation.game.game.score\[5\] _2324_ _2319_ vssd1 vssd1 vccd1 vccd1 _2336_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9201_ _0139_ _0411_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_7393_ net240 _2409_ _3016_ net433 net203 vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__o32a_1
XFILLER_0_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6344_ _2247_ _2250_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__nand2_1
X_9132_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[26\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9063_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[9\] net190 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[9\] sky130_fd_sc_hd__dfrtp_1
X_6275_ allocation.game.controller.drawBlock.counter\[4\] _2199_ vssd1 vssd1 vccd1
+ vccd1 _2200_ sky130_fd_sc_hd__xor2_1
X_5226_ _1148_ _1149_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nor2_1
X_8014_ net274 _3487_ _3523_ vssd1 vssd1 vccd1 vccd1 _3524_ sky130_fd_sc_hd__o21ai_1
X_5157_ _1077_ _1079_ _1080_ _0836_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__o211a_1
X_5088_ _0933_ _0935_ _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8916_ _4364_ _4365_ vssd1 vssd1 vccd1 vccd1 _4366_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8847_ _4295_ _4296_ vssd1 vssd1 vccd1 vccd1 _4297_ sky130_fd_sc_hd__and2b_1
X_8778_ net128 _3770_ _4225_ vssd1 vssd1 vccd1 vccd1 _4228_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7729_ net96 net66 vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__nand2_1
XANTENNA__7209__A _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8031__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8982__B _3219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9360__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7553__S net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7102__A1 allocation.game.controller.drawBlock.y_end\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7102__B2 allocation.game.controller.drawBlock.y_start\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6060_ net87 _0894_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__and2_1
X_5011_ _0924_ _0934_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__and2_1
X_6962_ _2712_ net91 _2711_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__and3b_1
XANTENNA__5102__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6893_ allocation.game.cactusDist.clock_div_inst0.counter\[3\] allocation.game.cactusDist.clock_div_inst0.counter\[2\]
+ allocation.game.cactusDist.clock_div_inst0.counter\[5\] allocation.game.cactusDist.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__or4_1
X_8701_ _0674_ _4151_ vssd1 vssd1 vccd1 vccd1 _4152_ sky130_fd_sc_hd__nand2_1
X_5913_ _1818_ _1820_ _1774_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__a21oi_1
X_5844_ _0723_ _0888_ _1768_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__or3b_1
X_8632_ _4072_ _4082_ vssd1 vssd1 vccd1 vccd1 _4083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8413__A _3256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8563_ net68 _3676_ vssd1 vssd1 vccd1 vccd1 _4014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4660__B allocation.game.controller.drawBlock.y_end\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8132__B net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7514_ _3073_ _3125_ _3058_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__or3b_1
X_5775_ _1634_ _1647_ _1646_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4726_ net229 allocation.game.cactusMove.x_dist\[2\] net227 vssd1 vssd1 vccd1 vccd1
+ _0653_ sky130_fd_sc_hd__a21oi_1
XANTENNA__8669__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8494_ _3903_ _3946_ net235 net233 net281 vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_47_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4657_ allocation.game.controller.drawBlock.y_start\[2\] allocation.game.controller.drawBlock.y_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7445_ net253 _3021_ allocation.game.lcdOutput.tft.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _3062_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7376_ allocation.game.cactusDist.lfsr1\[1\] allocation.game.cactusDist.lfsr2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4588_ _4456_ allocation.game.controller.v\[0\] vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__or2_1
X_6327_ _2250_ vssd1 vssd1 vccd1 vccd1 _2251_ sky130_fd_sc_hd__inv_2
X_9115_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[9\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9046_ clknet_leaf_3_clk allocation.game.dinoJump.next_dinoY\[0\] net195 vssd1 vssd1
+ vccd1 vccd1 allocation.game.collision.dinoY\[0\] sky130_fd_sc_hd__dfstp_2
X_6258_ _2108_ _2109_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8841__B2 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4675__X _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5209_ _0838_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__and2_1
X_6189_ _2112_ _2113_ _1810_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__a21o_1
XANTENNA__4835__B net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9233__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9383__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4570__B allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8832__B2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _1481_ _1484_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__and2b_1
X_4511_ allocation.game.bcd_ones\[3\] vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5491_ _1367_ _1369_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__xnor2_1
Xhold105 allocation.game.controller.init_module.delay_counter\[15\] vssd1 vssd1 vccd1
+ vccd1 net428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7230_ allocation.game.dinoJump.count\[16\] allocation.game.dinoJump.count\[17\]
+ _2901_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9106__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold116 allocation.game.cactusDist.clock_div_inst1.clk1 vssd1 vssd1 vccd1 vccd1 net439
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 allocation.game.controller.state\[5\] vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold127 allocation.game.cactus1size.clock_div_inst0.counter\[6\] vssd1 vssd1 vccd1
+ vccd1 net450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 allocation.game.cactus1size.clock_div_inst1.counter\[9\] vssd1 vssd1 vccd1
+ vccd1 net472 sky130_fd_sc_hd__dlygate4sd3_1
X_7161_ _2850_ _2855_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__nand2_1
X_7092_ allocation.game.controller.drawBlock.x_end\[4\] _2777_ _2779_ allocation.game.controller.drawBlock.y_end\[4\]
+ _0417_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6112_ _2007_ _2034_ _2033_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__a21o_1
XANTENNA__4936__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6834__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9256__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6043_ _1925_ _1966_ _1965_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7994_ net134 _3504_ vssd1 vssd1 vccd1 vccd1 _3505_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6945_ allocation.game.scoreCounter.clock_div.counter\[4\] allocation.game.scoreCounter.clock_div.counter\[3\]
+ _2396_ allocation.game.scoreCounter.clock_div.counter\[5\] vssd1 vssd1 vccd1 vccd1
+ _2702_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8339__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6876_ allocation.game.cactusDist.clock_div_inst1.counter\[7\] _2656_ _2658_ vssd1
+ vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5827_ _1748_ _1750_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__xnor2_1
X_8615_ net119 _4063_ _4065_ net97 vssd1 vssd1 vccd1 vccd1 _4066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8546_ net217 net115 vssd1 vssd1 vccd1 vccd1 _3997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5758_ _1682_ _1681_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_20_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4709_ net229 net227 allocation.game.cactusMove.x_dist\[2\] vssd1 vssd1 vccd1 vccd1
+ _0636_ sky130_fd_sc_hd__and3_1
X_8477_ net115 net51 _3881_ vssd1 vssd1 vccd1 vccd1 _3930_ sky130_fd_sc_hd__or3_1
X_5689_ net63 _1572_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__xnor2_1
X_7428_ net253 net252 vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7359_ allocation.game.lcdOutput.tft.remainingDelayTicks\[22\] _2998_ vssd1 vssd1
+ vccd1 vccd1 _2999_ sky130_fd_sc_hd__nor2_1
XANTENNA__4846__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9029_ clknet_leaf_4_clk _0154_ net187 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8027__C1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4565__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4603__A2 _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8053__A _4459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8988__A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9129__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9279__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _0901_ _0911_ _0915_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__a21oi_1
X_6730_ _2561_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6661_ net229 _2515_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_pixel\[2\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8400_ allocation.game.controller.v\[5\] net85 _3855_ vssd1 vssd1 vccd1 vccd1 _0386_
+ sky130_fd_sc_hd__a21o_1
X_6592_ net452 _2470_ net149 vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__o21ai_1
X_5612_ _0810_ _1536_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9380_ clknet_leaf_3_clk _0290_ net199 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight2\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_14_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8331_ net266 _3782_ vssd1 vssd1 vccd1 vccd1 _3795_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5543_ _1437_ _1465_ _1467_ _1409_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__o211a_1
XANTENNA__8410__B net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7847__A2 _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8262_ _2997_ _3733_ net55 vssd1 vssd1 vccd1 vccd1 _3734_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5474_ _1397_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__and2b_1
X_7213_ net84 _2892_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__and2_1
X_8193_ _0623_ _3683_ net113 vssd1 vssd1 vccd1 vccd1 _3684_ sky130_fd_sc_hd__a21oi_1
X_7144_ _2840_ _2846_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__or2_1
X_7075_ _2763_ _2778_ _2775_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__o21ai_1
X_6026_ _1948_ _1949_ _1950_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_1_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7977_ _0493_ _0500_ _3470_ vssd1 vssd1 vccd1 vccd1 _3489_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_25_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ allocation.game.cactusDist.clock_div_inst0.counter\[10\] _2690_ allocation.game.cactusDist.clock_div_inst0.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout55 _3000_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_2
XFILLER_0_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6859_ allocation.game.cactusDist.clock_div_inst1.counter\[1\] allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__nand2_1
Xfanout44 _3266_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_4
Xfanout88 _0759_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_2
Xfanout77 _2405_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_4
Xfanout99 _3190_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_4
Xfanout66 net67 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9421__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8529_ _3289_ _3305_ _3324_ net114 vssd1 vssd1 vccd1 vccd1 _3981_ sky130_fd_sc_hd__o31a_1
XFILLER_0_27_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7774__A1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload14 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload14/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7561__S net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5190_ net62 _1054_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__nor2_1
X_7900_ allocation.game.controller.drawBlock.counter\[10\] _3430_ vssd1 vssd1 vccd1
+ vccd1 _3432_ sky130_fd_sc_hd__nand2_1
X_8880_ _4305_ _4329_ _4310_ vssd1 vssd1 vccd1 vccd1 _4330_ sky130_fd_sc_hd__a21o_1
XANTENNA__9100__RESET_B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7831_ _2348_ _2358_ _2338_ vssd1 vssd1 vccd1 vccd1 _3389_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4974_ _0698_ _0898_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__and2_1
X_7762_ net66 net56 vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_19_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9501_ net286 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
X_6713_ net472 _2548_ net152 vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__o21ai_1
X_7693_ _3242_ _3243_ _3244_ _3247_ vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9444__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9432_ clknet_leaf_10_clk _0341_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6644_ allocation.game.cactusMove.count\[25\] allocation.game.cactusMove.count\[24\]
+ _2501_ allocation.game.cactusMove.count\[26\] vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8421__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_16
X_6575_ net145 _2461_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__nor2_2
X_9363_ clknet_leaf_5_clk _0012_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.bcd_tens\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8314_ _0488_ _3533_ _3778_ vssd1 vssd1 vccd1 vccd1 _3779_ sky130_fd_sc_hd__o21a_1
XANTENNA__7037__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5526_ _1450_ _1449_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__and2b_1
X_9294_ clknet_leaf_21_clk _0076_ net189 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5457_ _0754_ _0821_ _1379_ _1381_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__o2bb2ai_1
X_8245_ _2991_ _3722_ net54 vssd1 vssd1 vccd1 vccd1 _3723_ sky130_fd_sc_hd__a21o_1
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_4
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
Xfanout223 allocation.game.cactusMove.pixel\[6\] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
X_8176_ _0652_ net77 _3668_ _0683_ vssd1 vssd1 vccd1 vccd1 _3669_ sky130_fd_sc_hd__o22a_1
XANTENNA__5700__B1 _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5388_ _1293_ _1295_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout256 allocation.game.lcdOutput.tft.spiDataSet vssd1 vssd1 vccd1 vccd1 net256
+ sky130_fd_sc_hd__clkbuf_4
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
X_7127_ _2832_ _2833_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__nor2_1
Xfanout245 allocation.game.lcdOutput.tft.initSeqCounter\[5\] vssd1 vssd1 vccd1 vccd1
+ net245 sky130_fd_sc_hd__buf_2
X_7058_ _0443_ allocation.game.controller.drawBlock.idx\[1\] allocation.game.controller.drawBlock.idx\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__or3_2
Xfanout278 allocation.game.collision.dinoY\[1\] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
Xfanout267 allocation.game.collision.dinoY\[5\] vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
X_6009_ _1927_ _1932_ _1933_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5939__B _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9520__305 vssd1 vssd1 vccd1 vccd1 _9520__305/HI net305 sky130_fd_sc_hd__conb_1
XFILLER_0_33_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8331__A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4990__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9317__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7556__S net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4690_ net222 _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6360_ net277 _2282_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__or2_1
X_5311_ _1017_ _1026_ _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8030_ net266 _3521_ vssd1 vssd1 vccd1 vccd1 _3539_ sky130_fd_sc_hd__nor2_1
X_6291_ _2190_ _2191_ _2193_ allocation.game.controller.drawBlock.counter\[7\] _2215_
+ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__o221a_1
XANTENNA__8475__A2 _3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5242_ _1160_ _1164_ _1165_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5173_ net60 _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5105__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 en vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8932_ _4331_ _4351_ _4381_ vssd1 vssd1 vccd1 vccd1 _4382_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5759__B _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8863_ _0467_ net35 _3811_ _4305_ _4312_ vssd1 vssd1 vccd1 vccd1 _4313_ sky130_fd_sc_hd__o311a_1
XFILLER_0_17_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7814_ net234 allocation.game.bcd_ones\[0\] net232 vssd1 vssd1 vccd1 vccd1 _3375_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8794_ net261 _3540_ vssd1 vssd1 vccd1 vccd1 _4244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4957_ _0863_ _0881_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7745_ net114 _3304_ _3305_ _3306_ vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8163__B2 allocation.game.controller.drawBlock.x_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4888_ _0811_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__nand2_2
X_7676_ allocation.game.lcdOutput.framebufferIndex\[6\] net48 vssd1 vssd1 vccd1 vccd1
+ _3238_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9415_ clknet_leaf_13_clk _0324_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.idx\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6627_ allocation.game.cactusMove.count\[19\] _2492_ _2494_ vssd1 vssd1 vccd1 vccd1
+ allocation.game.cactusMove.n_count\[19\] sky130_fd_sc_hd__o21a_1
XFILLER_0_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7990__A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9346_ clknet_leaf_5_clk _0278_ net173 vssd1 vssd1 vccd1 vccd1 allocation.game.game.score\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_6558_ _2447_ _2415_ _2446_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[18\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6489_ allocation.game.scoreCounter.clock_div.counter\[24\] allocation.game.scoreCounter.clock_div.counter\[23\]
+ _2403_ allocation.game.scoreCounter.clock_div.counter\[25\] vssd1 vssd1 vccd1 vccd1
+ _2404_ sky130_fd_sc_hd__a31oi_1
X_9277_ clknet_leaf_2_clk _0265_ net181 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.lfsr2\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_5509_ _1433_ _1432_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__and2b_1
XANTENNA__4838__B _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8228_ allocation.game.lcdOutput.tft.remainingDelayTicks\[6\] _2986_ vssd1 vssd1
+ vccd1 vccd1 _3712_ sky130_fd_sc_hd__nand2_1
X_8159_ allocation.game.controller.state\[1\] _3648_ _3649_ _3656_ vssd1 vssd1 vccd1
+ vccd1 _3657_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4854__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8926__B1 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8061__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4748__B net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5860_ _0800_ _0899_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__nor2_1
X_4811_ _0555_ _0568_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5791_ _1662_ _1715_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4742_ _0664_ _0668_ net217 vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__o21ai_2
X_7530_ _3060_ _3137_ _3139_ _3133_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__a211o_1
X_4673_ allocation.game.controller.drawBlock.y_end\[7\] allocation.game.controller.drawBlock.y_start\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7461_ _4463_ net252 vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__nor2_1
X_6412_ allocation.game.game.score\[5\] _2331_ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9200_ _0138_ _0410_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__8696__A2 _3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7392_ net243 net239 _2413_ net204 vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__o31ai_1
X_6343_ net259 net263 vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__nand2_1
X_9131_ clknet_leaf_2_clk allocation.game.cactusMove.n_count\[25\] net177 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[25\] sky130_fd_sc_hd__dfrtp_1
X_9062_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[8\] net190 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6274_ _2085_ _2095_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__nand2_1
X_5225_ _1148_ _1149_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__and2_1
X_8013_ _3521_ _3522_ vssd1 vssd1 vccd1 vccd1 _3523_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5156_ _0836_ _1080_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5087_ _0973_ _1010_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__xnor2_1
X_8915_ net264 _4352_ net261 vssd1 vssd1 vccd1 vccd1 _4365_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4961__X _0886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8846_ net133 _4457_ vssd1 vssd1 vccd1 vccd1 _4296_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4680__Y allocation.game.cactus1size.clock_div_inst0.reset vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_5989_ _1866_ _1868_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__xnor2_1
X_8777_ _4226_ vssd1 vssd1 vccd1 vccd1 _4227_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7728_ net117 _3288_ vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7659_ _3217_ _3214_ _3212_ vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__mux2_1
X_9329_ clknet_leaf_6_clk _0112_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__7225__A _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8056__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4658__A_N allocation.game.controller.drawBlock.y_end\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4871__X _0796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9526__311 vssd1 vssd1 vccd1 vccd1 _9526__311/HI net311 sky130_fd_sc_hd__conb_1
XANTENNA__8375__B2 allocation.game.controller.drawBlock.y_end\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5189__A1 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5010_ _0924_ _0934_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nor2_1
XANTENNA__9035__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6961_ allocation.game.scoreCounter.clock_div.counter\[11\] allocation.game.scoreCounter.clock_div.counter\[10\]
+ _2708_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__and3_1
X_8700_ net112 _3670_ vssd1 vssd1 vccd1 vccd1 _4151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8366__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6892_ net333 _2666_ _2668_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__a21oi_1
X_5912_ _0896_ _1834_ _1835_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__nand3_2
X_8631_ net225 _2519_ vssd1 vssd1 vccd1 vccd1 _4082_ sky130_fd_sc_hd__or2_1
X_5843_ _0715_ _0886_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8562_ _4011_ _4012_ vssd1 vssd1 vccd1 vccd1 _4013_ sky130_fd_sc_hd__or2_1
X_5774_ _1683_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__or2_1
X_7513_ net248 _3046_ _3042_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__o21a_1
XANTENNA__6129__B1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4725_ _0635_ _0646_ _0647_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o21a_1
X_8493_ _3360_ _3938_ _3945_ _3926_ _3933_ vssd1 vssd1 vccd1 vccd1 _3946_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4656_ allocation.game.controller.drawBlock.y_start\[3\] allocation.game.controller.drawBlock.y_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout215_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7444_ net253 net248 vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__or2_1
X_4587_ net280 _0519_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nand2_1
X_7375_ allocation.game.lcdOutput.tft.remainingDelayTicks\[22\] _2998_ net329 vssd1
+ vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9114_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[8\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[8\] sky130_fd_sc_hd__dfrtp_1
X_6326_ net265 _2243_ _2249_ net271 vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9045_ clknet_leaf_7_clk _0170_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_6257_ allocation.game.controller.drawBlock.counter\[13\] _2181_ vssd1 vssd1 vccd1
+ vccd1 _2182_ sky130_fd_sc_hd__nand2_1
X_5208_ _0780_ _0784_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__xnor2_1
X_6188_ _1807_ _1809_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__xnor2_1
X_5139_ _0809_ _0822_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__and2_1
XANTENNA__5947__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8829_ net258 _4278_ vssd1 vssd1 vccd1 vccd1 _4279_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7096__A1 allocation.game.controller.drawBlock.y_end\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7402__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9058__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5490_ _1414_ _1412_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__and2b_1
X_4510_ allocation.game.bcd_ones\[0\] vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
Xhold106 allocation.game.controller.drawBlock.y_end\[0\] vssd1 vssd1 vccd1 vccd1 net429
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 allocation.game.cactusDist.clock_div_inst0.counter\[12\] vssd1 vssd1 vccd1
+ vccd1 net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 allocation.game.controller.drawBlock.x_start\[3\] vssd1 vssd1 vccd1 vccd1
+ net451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 allocation.game.cactusHeight2\[4\] vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7160_ _2847_ _2858_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6111_ _0769_ _0894_ _1961_ _1960_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__a31o_1
X_7091_ allocation.game.controller.drawBlock.x_start\[4\] _2772_ _2787_ allocation.game.controller.drawBlock.y_start\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6042_ _1925_ _1965_ _1966_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__nor3_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7993_ _0490_ _0499_ vssd1 vssd1 vccd1 vccd1 _3504_ sky130_fd_sc_hd__nor2_1
XANTENNA__8051__A3 _3559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8339__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6944_ net372 _2397_ _2701_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6875_ allocation.game.cactusDist.clock_div_inst1.counter\[7\] _2656_ net159 vssd1
+ vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__a21oi_1
X_8614_ _2524_ _4064_ vssd1 vssd1 vccd1 vccd1 _4065_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5826_ _1750_ _1748_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__and2b_1
X_5757_ _1630_ _1631_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8545_ _2861_ _3995_ _3342_ vssd1 vssd1 vccd1 vccd1 _3996_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4708_ net226 allocation.game.cactusMove.x_dist\[4\] vssd1 vssd1 vccd1 vccd1 _0635_
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout120_X net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8476_ _3297_ _3880_ _3883_ vssd1 vssd1 vccd1 vccd1 _3929_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5688_ net63 _1612_ _1611_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__a21bo_1
X_7427_ _0430_ _3042_ _0429_ net245 vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__o211a_1
X_4639_ _0554_ _0568_ _0553_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7358_ allocation.game.lcdOutput.tft.remainingDelayTicks\[21\] _2997_ vssd1 vssd1
+ vccd1 vccd1 _2998_ sky130_fd_sc_hd__or2_1
X_7289_ _2947_ _2948_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__nor2_1
X_6309_ _2156_ _2233_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__nor2_2
XANTENNA__8275__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9028_ clknet_leaf_4_clk _0153_ net185 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout78_A _0796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9350__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8750__A1 _3228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7384__S _2973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7559__S net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4990_ net124 net102 _0913_ net78 vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__a31o_1
X_6660_ net151 _2461_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6591_ allocation.game.cactusMove.count\[5\] allocation.game.cactusMove.count\[6\]
+ _2468_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__and3_1
X_5611_ _1496_ _1498_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8330_ _3792_ _3793_ vssd1 vssd1 vccd1 vccd1 _3794_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5542_ _1406_ _1408_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9223__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8261_ allocation.game.lcdOutput.tft.remainingDelayTicks\[19\] _2995_ allocation.game.lcdOutput.tft.remainingDelayTicks\[20\]
+ vssd1 vssd1 vccd1 vccd1 _3733_ sky130_fd_sc_hd__o21ai_1
X_5473_ _1347_ _1349_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__xnor2_1
X_7212_ allocation.game.dinoJump.count\[9\] allocation.game.dinoJump.count\[10\] allocation.game.dinoJump.count\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__and3_1
X_8192_ net222 _0621_ vssd1 vssd1 vccd1 vccd1 _3683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7143_ allocation.game.lcdOutput.framebufferIndex\[12\] _2839_ allocation.game.lcdOutput.framebufferIndex\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__a21oi_1
X_7074_ allocation.game.controller.color\[10\] _2786_ _2792_ allocation.game.controller.color\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__a22o_1
XANTENNA__9373__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6025_ _0716_ _0905_ _0907_ net110 vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7976_ net277 _3473_ net134 vssd1 vssd1 vccd1 vccd1 _3488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ allocation.game.cactusDist.clock_div_inst0.counter\[10\] _2690_ _2692_ vssd1
+ vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9047__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout56 net57 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout45 _3266_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_2
X_6858_ allocation.game.cactusDist.clock_div_inst1.counter\[0\] net152 _2646_ vssd1
+ vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__and3b_1
Xfanout34 _3272_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_2
Xfanout78 _0796_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_4
X_5809_ _0769_ _0907_ _1732_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__a21o_1
Xfanout67 _3209_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_2
XFILLER_0_18_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout89 _0671_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8528_ _3339_ _3979_ _3958_ vssd1 vssd1 vccd1 vccd1 _3980_ sky130_fd_sc_hd__a21oi_1
X_6789_ allocation.game.cactus2size.clock_div_inst1.counter\[6\] _2600_ vssd1 vssd1
+ vccd1 vccd1 _2601_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8459_ _3324_ _3892_ vssd1 vssd1 vccd1 vccd1 _3912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4592__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9246__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload15 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_16
XANTENNA__9396__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7830_ _2348_ _2358_ vssd1 vssd1 vccd1 vccd1 _3388_ sky130_fd_sc_hd__and2_1
X_4973_ _0592_ _0696_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__nand2_1
X_7761_ _3288_ _3320_ _3321_ net118 vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9500_ net285 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
X_7692_ allocation.game.lcdOutput.framebufferIndex\[4\] _3239_ _3251_ _3253_ vssd1
+ vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__and4_1
X_6712_ allocation.game.cactus1size.clock_div_inst1.counter\[9\] _2548_ vssd1 vssd1
+ vccd1 vccd1 _2549_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9431_ clknet_leaf_10_clk _0340_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_6643_ allocation.game.cactusMove.count\[25\] _2502_ _2504_ vssd1 vssd1 vccd1 vccd1
+ allocation.game.cactusMove.n_count\[25\] sky130_fd_sc_hd__o21a_1
XFILLER_0_15_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8714__A1 net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload9 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_16
XFILLER_0_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9362_ clknet_leaf_12_clk _0011_ net204 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6574_ _2453_ _2454_ _2455_ _2460_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__nor4_4
XFILLER_0_14_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout128_A allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_8313_ _0488_ _0504_ vssd1 vssd1 vccd1 vccd1 _3778_ sky130_fd_sc_hd__nand2_1
X_5525_ _0838_ _1444_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9293_ clknet_leaf_2_clk _0267_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.clk1
+ sky130_fd_sc_hd__dfxtp_1
X_5456_ _0865_ _1380_ _0866_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__a21o_1
X_8244_ allocation.game.lcdOutput.tft.remainingDelayTicks\[12\] _2990_ vssd1 vssd1
+ vccd1 vccd1 _3722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout202 net216 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5700__B2 _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5700__A1 _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8149__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8175_ net164 _0687_ _3667_ vssd1 vssd1 vccd1 vccd1 _3668_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5387_ _1310_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__or2_1
Xfanout224 allocation.game.cactusMove.pixel\[5\] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
X_7126_ allocation.game.lcdOutput.framebufferIndex\[6\] _2830_ vssd1 vssd1 vccd1 vccd1
+ _2833_ sky130_fd_sc_hd__nor2_1
Xfanout246 allocation.game.lcdOutput.tft.initSeqCounter\[5\] vssd1 vssd1 vccd1 vccd1
+ net246 sky130_fd_sc_hd__clkbuf_2
Xfanout235 allocation.game.cactus1size.state\[0\] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
X_7057_ _2771_ _2773_ vssd1 vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__nor2_2
Xfanout279 allocation.game.collision.dinoY\[1\] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout257 allocation.game.cactusMove.x_dist\[1\] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input2_A gpio_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 net271 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
XANTENNA__9119__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6008_ _1890_ _1931_ _1930_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5301__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8953__A1 _3208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7959_ net280 net278 vssd1 vssd1 vccd1 vccd1 _3472_ sky130_fd_sc_hd__or2_1
XANTENNA__9269__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8705__B2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8705__A1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5211__A _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5310_ _1233_ _1234_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6290_ allocation.game.controller.drawBlock.counter\[7\] _2193_ _2195_ allocation.game.controller.drawBlock.counter\[6\]
+ _2214_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_12_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5241_ _1160_ _1164_ _1165_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__a21oi_1
X_5172_ _1068_ _1087_ _1089_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_3_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 gpio_in[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8931_ _4371_ _4379_ _4380_ vssd1 vssd1 vccd1 vccd1 _4381_ sky130_fd_sc_hd__nand3_1
XANTENNA__9411__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7199__B1 _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8862_ net270 net43 _4306_ _4307_ _4311_ vssd1 vssd1 vccd1 vccd1 _4312_ sky130_fd_sc_hd__o221a_1
X_8793_ _4242_ vssd1 vssd1 vccd1 vccd1 _4243_ sky130_fd_sc_hd__inv_2
X_7813_ net235 net233 net199 _3374_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__and4_1
X_7744_ net114 _3289_ _3291_ vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4956_ _0826_ _0879_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4887_ _0809_ _0810_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__nand2b_1
X_7675_ net48 vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__inv_2
X_9414_ clknet_leaf_13_clk _0323_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.idx\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_6626_ allocation.game.cactusMove.count\[19\] _2492_ net145 vssd1 vssd1 vccd1 vccd1
+ _2494_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9345_ clknet_leaf_5_clk _0277_ net173 vssd1 vssd1 vccd1 vccd1 allocation.game.game.score\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_6557_ allocation.game.dinoJump.dinoDelay\[17\] allocation.game.dinoJump.dinoDelay\[18\]
+ _2443_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5508_ _1379_ _1381_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__xnor2_1
X_6488_ _2399_ _2402_ _2395_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9276_ clknet_leaf_2_clk _0264_ net181 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.lfsr2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_5439_ _1312_ _1314_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__and2_1
X_8227_ _0420_ _3001_ _3033_ _3711_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__o211a_1
X_8158_ allocation.game.controller.state\[2\] _3652_ _3653_ _3655_ vssd1 vssd1 vccd1
+ vccd1 _3656_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7109_ allocation.game.controller.init_module.idx\[0\] _0425_ _2757_ vssd1 vssd1
+ vccd1 vccd1 _2821_ sky130_fd_sc_hd__or3_2
X_8089_ _3591_ _3592_ allocation.game.controller.drawBlock.x_end\[1\] net206 vssd1
+ vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__9409__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9091__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4854__B _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6165__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9434__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7968__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ _0720_ _0734_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5790_ net63 _1661_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4741_ _0665_ _0667_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__and2b_1
X_4672_ _0578_ _0601_ _0577_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a21o_2
XFILLER_0_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7460_ _3052_ _3075_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__nand2_1
X_6411_ _2333_ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7391_ net385 net206 _3015_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9130_ clknet_leaf_2_clk allocation.game.cactusMove.n_count\[24\] net181 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6342_ _2263_ _2265_ _2252_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9061_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[7\] net192 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[7\] sky130_fd_sc_hd__dfrtp_1
X_6273_ allocation.game.controller.drawBlock.counter\[5\] _2197_ vssd1 vssd1 vccd1
+ vccd1 _2198_ sky130_fd_sc_hd__xnor2_1
X_5224_ _1076_ _1090_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__xnor2_1
X_8012_ net273 net269 vssd1 vssd1 vccd1 vccd1 _3522_ sky130_fd_sc_hd__or2_2
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout195_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5155_ _0834_ _0835_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8081__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5086_ _1010_ _0973_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__and2b_1
X_8914_ _0467_ _4352_ vssd1 vssd1 vccd1 vccd1 _4364_ sky130_fd_sc_hd__and2_1
X_8845_ net133 _4457_ vssd1 vssd1 vccd1 vccd1 _4295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _1909_ _1912_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout150_X net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8776_ _3770_ _4225_ net128 vssd1 vssd1 vccd1 vccd1 _4226_ sky130_fd_sc_hd__a21oi_1
X_4939_ _0806_ _0813_ _0811_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_30_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7727_ net96 net74 vssd1 vssd1 vccd1 vccd1 _3289_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_44_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9307__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7658_ allocation.game.lcdOutput.framebufferIndex\[8\] net56 vssd1 vssd1 vccd1 vccd1
+ _3220_ sky130_fd_sc_hd__and2_1
X_6609_ _2482_ _2483_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[12\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7589_ allocation.game.cactus2size.clock_div_inst1.clk1 allocation.game.cactus2size.lfsr2\[1\]
+ allocation.game.cactus2size.lfsr2\[0\] vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__a21oi_1
X_9328_ clknet_leaf_6_clk _0111_ net174 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9259_ clknet_leaf_2_clk _0261_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.clk1
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__A _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout63_X net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8800__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6320__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6960_ allocation.game.scoreCounter.clock_div.counter\[11\] _2710_ vssd1 vssd1 vccd1
+ vccd1 _2711_ sky130_fd_sc_hd__or2_1
X_5911_ _1834_ _1835_ _0896_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__a21o_1
XANTENNA__4781__Y _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6891_ net333 _2666_ net152 vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__o21ai_1
XANTENNA__6377__A1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6377__B2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8630_ _2519_ _4061_ vssd1 vssd1 vccd1 vccd1 _4081_ sky130_fd_sc_hd__xnor2_1
X_5842_ _1723_ _1724_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8561_ net56 _3608_ vssd1 vssd1 vccd1 vccd1 _4012_ sky130_fd_sc_hd__nor2_1
X_5773_ _1696_ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__and2_1
XANTENNA__6129__A1 _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4724_ _0649_ _0650_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__or2_1
X_7512_ _3120_ _3121_ _3123_ vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__a21o_1
XANTENNA__6129__B2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8492_ _3909_ _3944_ vssd1 vssd1 vccd1 vccd1 _3945_ sky130_fd_sc_hd__nand2b_1
X_4655_ _0583_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__nand2b_2
X_7443_ net247 net246 vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__nor2_2
X_4586_ net233 _0521_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoY\[2\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout110_A _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7374_ _2999_ _3007_ _3001_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout208_A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9113_ clknet_leaf_7_clk allocation.game.cactusMove.n_count\[7\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[7\] sky130_fd_sc_hd__dfrtp_1
X_6325_ _2239_ _2248_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9044_ clknet_leaf_7_clk _0169_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6256_ _1905_ _2110_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5207_ _0784_ _0780_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__and2b_1
X_6187_ _1857_ _2111_ _1856_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__a21o_1
X_5138_ _1061_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__nor2_1
X_5069_ _0989_ _0992_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__and2_1
XANTENNA__8357__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8828_ _0468_ _4277_ vssd1 vssd1 vccd1 vccd1 _4278_ sky130_fd_sc_hd__nor2_1
X_8759_ _3305_ _3882_ vssd1 vssd1 vccd1 vccd1 _4209_ sky130_fd_sc_hd__and2_1
XANTENNA__8109__A2 _3609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 allocation.game.cactus2size.clock_div_inst1.counter\[3\] vssd1 vssd1 vccd1
+ vccd1 net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 allocation.game.cactusMove.count\[6\] vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 allocation.game.cactus1size.clock_div_inst1.counter\[6\] vssd1 vssd1 vccd1
+ vccd1 net441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6110_ _2007_ _2033_ _2034_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__nand3_1
X_7090_ _2802_ _2805_ _2806_ _2801_ vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__o31a_1
X_6041_ _1922_ _1923_ _1924_ _1863_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9152__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7992_ _0487_ _0489_ _0499_ vssd1 vssd1 vccd1 vccd1 _3503_ sky130_fd_sc_hd__and3_1
X_6943_ allocation.game.scoreCounter.clock_div.counter\[4\] _2397_ net91 vssd1 vssd1
+ vccd1 vccd1 _2701_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6225__A _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6874_ _2656_ _2657_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8613_ net220 _2375_ vssd1 vssd1 vccd1 vccd1 _4064_ sky130_fd_sc_hd__nor2_1
X_5825_ _1698_ _1749_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5756_ _0990_ _1668_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__o21ai_1
X_8544_ net132 net130 net126 net44 net41 vssd1 vssd1 vccd1 vccd1 _3995_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_20_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7327__Y _2973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4707_ _0632_ _0633_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5687_ _1609_ _1610_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__xnor2_1
X_8475_ _3285_ _3362_ _3909_ vssd1 vssd1 vccd1 vccd1 _3928_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_20_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4638_ _0557_ _0567_ _0556_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__a21o_1
X_7426_ _0430_ _3042_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__nor2_1
XANTENNA__4648__A_N allocation.game.controller.drawBlock.y_end\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ _0486_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nand2_1
X_7357_ allocation.game.lcdOutput.tft.remainingDelayTicks\[20\] _2996_ vssd1 vssd1
+ vccd1 vccd1 _2997_ sky130_fd_sc_hd__or2_1
X_7288_ allocation.game.controller.init_module.delay_counter\[10\] _2946_ net122 vssd1
+ vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__o21ai_1
X_6308_ _2132_ _2159_ _2232_ _2157_ _2158_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__a2111o_1
XANTENNA__8275__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9027_ clknet_leaf_9_clk _0152_ net185 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6239_ _2125_ _2126_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__nor2_1
XANTENNA__8027__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9025__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9175__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7241__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6590_ _2470_ _2471_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5610_ _1065_ _1534_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5541_ _1465_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8260_ _3034_ _3732_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__or2_1
X_7211_ allocation.game.dinoJump.count\[11\] _2889_ _2891_ vssd1 vssd1 vccd1 vccd1
+ _2892_ sky130_fd_sc_hd__o21ba_1
X_5472_ _0864_ _1391_ _1396_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8191_ _0663_ _3681_ _0682_ vssd1 vssd1 vccd1 vccd1 _3682_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4947__B _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7142_ _2842_ _2844_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkload12_A clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7073_ _2778_ _2785_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__nor2_1
X_6024_ _0741_ _0904_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__nor2_1
X_9511__296 vssd1 vssd1 vccd1 vccd1 _9511__296/HI net296 sky130_fd_sc_hd__conb_1
X_7975_ net277 _3473_ vssd1 vssd1 vccd1 vccd1 _3487_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ allocation.game.cactusDist.clock_div_inst0.counter\[10\] _2690_ net160 vssd1
+ vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout46 _3256_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_4
Xfanout35 net36 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_18_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6857_ _2646_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout79 _0796_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_2
X_5808_ _0770_ _0908_ _1732_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__or3b_1
Xfanout57 _3219_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_4
Xfanout68 net69 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_4
X_6788_ net162 _2599_ _2600_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__nor3_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9048__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5739_ net63 _1612_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__xnor2_1
X_8527_ _3288_ _3978_ _3905_ net117 vssd1 vssd1 vccd1 vccd1 _3979_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8458_ _3869_ _3909_ _3910_ vssd1 vssd1 vccd1 vccd1 _3911_ sky130_fd_sc_hd__or3_1
X_8389_ allocation.game.controller.v\[2\] net84 _3847_ vssd1 vssd1 vccd1 vccd1 _0383_
+ sky130_fd_sc_hd__a21o_1
X_7409_ allocation.game.lcdOutput.tft.state\[2\] allocation.game.lcdOutput.tft.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__nor2_1
XANTENNA__4873__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8723__A2 net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload16/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7760_ net117 _3321_ vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_19_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4972_ _0896_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__inv_2
X_7691_ _3252_ vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__inv_2
X_6711_ net159 _2547_ _2548_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__nor3_1
X_9430_ clknet_leaf_11_clk _0339_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_6642_ allocation.game.cactusMove.count\[25\] _2502_ net145 vssd1 vssd1 vccd1 vccd1
+ _2504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9361_ clknet_leaf_12_clk _0010_ net201 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8312_ _3593_ _3766_ _3777_ net197 allocation.game.controller.drawBlock.y_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__o32a_1
X_6573_ _2456_ _2457_ _2458_ _2459_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9340__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5524_ _0778_ _0888_ _1445_ _1448_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9292_ clknet_leaf_0_clk _0094_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8478__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5455_ _0778_ _0797_ _0832_ _0843_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8243_ _3035_ _3721_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__nand2_1
X_8174_ _0643_ _0656_ vssd1 vssd1 vccd1 vccd1 _3667_ sky130_fd_sc_hd__nand2_1
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_4
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
XANTENNA__5700__A2 _0886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7125_ allocation.game.lcdOutput.framebufferIndex\[6\] _2830_ vssd1 vssd1 vccd1 vccd1
+ _2832_ sky130_fd_sc_hd__and2_1
X_5386_ _1303_ _1305_ _1309_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__nor3_1
Xfanout236 allocation.game.controller.drawBlock.init_done vssd1 vssd1 vccd1 vccd1
+ net236 sky130_fd_sc_hd__clkbuf_4
Xfanout225 allocation.game.cactusMove.pixel\[5\] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
Xfanout247 allocation.game.lcdOutput.tft.initSeqCounter\[4\] vssd1 vssd1 vccd1 vccd1
+ net247 sky130_fd_sc_hd__clkbuf_4
XANTENNA__9490__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout258 net260 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_4
X_7056_ allocation.game.controller.drawBlock.x_start\[0\] _2772_ _2775_ vssd1 vssd1
+ vccd1 vccd1 _2776_ sky130_fd_sc_hd__a21bo_1
Xfanout269 net271 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6007_ _1890_ _1930_ _1931_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7958_ _0496_ _0523_ net134 vssd1 vssd1 vccd1 vccd1 _3471_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7889_ _3423_ _3424_ allocation.game.controller.drawBlock.counter\[6\] net108 vssd1
+ vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a2bb2o_1
X_6909_ allocation.game.cactusDist.clock_div_inst0.counter\[3\] allocation.game.cactusDist.clock_div_inst0.counter\[4\]
+ _2678_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7913__B1 _3409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7244__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5455__A1 _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9213__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9363__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7380__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5240_ _1106_ _1108_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7683__A2 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5171_ _1094_ _1095_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8930_ _4216_ _4244_ _3875_ _4209_ _4215_ vssd1 vssd1 vccd1 vccd1 _4380_ sky130_fd_sc_hd__o2111a_1
Xinput3 gpio_in[1] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XANTENNA__5759__D _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8861_ net38 _4304_ _4309_ vssd1 vssd1 vccd1 vccd1 _4311_ sky130_fd_sc_hd__o21a_1
X_7812_ _3364_ _3368_ _3373_ _3354_ _3269_ vssd1 vssd1 vccd1 vccd1 _3374_ sky130_fd_sc_hd__a32o_1
X_8792_ _3521_ _3760_ vssd1 vssd1 vccd1 vccd1 _4242_ sky130_fd_sc_hd__and2_1
X_4955_ _0826_ _0879_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__nand2b_1
XANTENNA__4960__B _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7743_ net48 _3293_ net50 vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout238_A allocation.game.controller.block_done vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4886_ _0810_ _0809_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__nand2b_1
X_7674_ _3233_ _3235_ vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__or2_1
X_9413_ clknet_leaf_13_clk _0322_ net211 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.idx\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_6625_ _2492_ _2493_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[18\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9344_ clknet_leaf_4_clk _0276_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.game.score\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_6556_ allocation.game.dinoJump.dinoDelay\[17\] _2443_ allocation.game.dinoJump.dinoDelay\[18\]
+ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__a21o_1
X_5507_ _1430_ _1431_ _1427_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__a21o_1
X_9275_ clknet_leaf_4_clk _0263_ net187 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.lfsr1\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6487_ _2389_ _2401_ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__nor2_1
X_8226_ _2986_ _3710_ vssd1 vssd1 vccd1 vccd1 _3711_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5438_ _1343_ _1362_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__nand2_1
X_8157_ net239 _3654_ _3597_ allocation.game.controller.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _3655_ sky130_fd_sc_hd__a211o_1
X_5369_ _1232_ _1241_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__and2_1
X_7108_ _2818_ _2819_ allocation.game.controller.init_module.delay_counter\[17\] allocation.game.controller.init_module.delay_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__o211a_1
X_8088_ net113 net77 vssd1 vssd1 vccd1 vccd1 _3593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7039_ _0424_ _2759_ _2756_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__a21o_1
XANTENNA__6634__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9236__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9386__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5982__A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8862__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4740_ _0664_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4671_ _0581_ _0600_ _0580_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9109__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7390_ net203 net101 vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__nand2_1
X_6410_ _2319_ _2327_ _2331_ _2332_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__a22oi_2
XANTENNA__8550__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6341_ _2261_ _2264_ _2259_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9060_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[6\] net192 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6272_ _2097_ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__nand2_1
X_5223_ _1130_ _1147_ _1129_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a21bo_1
X_8011_ net272 net270 vssd1 vssd1 vccd1 vccd1 _3521_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9259__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5154_ _0846_ _1078_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout188_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5085_ _1007_ _1009_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8369__B1 _0541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8913_ net41 _4353_ _4354_ _4361_ _4362_ vssd1 vssd1 vccd1 vccd1 _4363_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8844_ net258 _4278_ _4290_ _4293_ vssd1 vssd1 vccd1 vccd1 _4294_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4971__A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5987_ _1909_ _1910_ _1911_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__nand3_1
X_8775_ net272 _3760_ vssd1 vssd1 vccd1 vccd1 _4225_ sky130_fd_sc_hd__nand2_1
X_4938_ _0861_ _0862_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__or2_1
X_7726_ net99 _3200_ vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__nor2_2
X_4869_ _0771_ _0777_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7657_ _3212_ _3214_ _3216_ vssd1 vssd1 vccd1 vccd1 _3219_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6608_ allocation.game.cactusMove.count\[12\] _2480_ net147 vssd1 vssd1 vccd1 vccd1
+ _2483_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7588_ net144 _3166_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9327_ clknet_leaf_6_clk _0110_ net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6539_ allocation.game.dinoJump.dinoDelay\[11\] _2432_ allocation.game.dinoJump.dinoDelay\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9258_ clknet_leaf_0_clk _0066_ net176 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8209_ _0680_ _3647_ _0683_ vssd1 vssd1 vccd1 vccd1 _3698_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9189_ clknet_leaf_15_clk _0251_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9401__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7099__B1 _0417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8835__B2 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8835__A1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9420__Q allocation.game.controller.drawBlock.y_start\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5910_ _1787_ _1833_ _1832_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__a21o_1
X_6890_ _2666_ _2667_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5841_ _1728_ _1729_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8560_ net58 _3609_ vssd1 vssd1 vccd1 vccd1 _4011_ sky130_fd_sc_hd__nor2_1
X_5772_ _1681_ _1682_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__xnor2_1
X_4723_ net112 _0648_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8491_ _3287_ _3332_ _3868_ _3943_ vssd1 vssd1 vccd1 vccd1 _3944_ sky130_fd_sc_hd__a31o_1
X_7511_ net245 _3049_ _3122_ allocation.game.lcdOutput.tft.initSeqCounter\[4\] vssd1
+ vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7442_ _3055_ _3056_ _3058_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__and3_1
X_4654_ allocation.game.controller.drawBlock.y_end\[4\] allocation.game.controller.drawBlock.y_start\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9081__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4585_ net106 _0518_ _0520_ net235 vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__o211a_1
X_7373_ allocation.game.lcdOutput.tft.remainingDelayTicks\[22\] _2998_ vssd1 vssd1
+ vccd1 vccd1 _3007_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9112_ clknet_leaf_7_clk allocation.game.cactusMove.n_count\[6\] net184 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4560__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout103_A _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6324_ allocation.game.cactusHeight2\[3\] _2238_ allocation.game.cactusHeight2\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__a21oi_1
X_9043_ clknet_leaf_7_clk _0168_ net183 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_6255_ _1857_ _2111_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5206_ _1129_ _1130_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__nand2_1
X_6186_ _1905_ _2110_ _1904_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__o21ai_1
X_5137_ _1051_ _1055_ _1060_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nor3_1
X_5068_ _0989_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8827_ net268 _3770_ vssd1 vssd1 vccd1 vccd1 _4277_ sky130_fd_sc_hd__nand2_1
X_8758_ _4208_ net199 net151 vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__and3b_1
XFILLER_0_30_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7709_ net37 _3264_ vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__nor2_2
XANTENNA__9424__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8689_ _4118_ _4137_ _4138_ vssd1 vssd1 vccd1 vccd1 _4140_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4876__A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8348__A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5500__A _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold108 allocation.game.controller.drawBlock.x_start\[5\] vssd1 vssd1 vccd1 vccd1
+ net431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 allocation.game.dinoJump.count\[16\] vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6040_ _1962_ _1964_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8545__X _3996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7991_ _3500_ _3501_ _3502_ net203 net400 vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__o32a_1
X_6942_ _2397_ net91 _2700_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__and3b_1
XANTENNA__6506__A _0464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6873_ net478 _2655_ net152 vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9447__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5824_ _1696_ _1697_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__nor2_1
X_8612_ net217 _2524_ vssd1 vssd1 vccd1 vccd1 _4063_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_33_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7337__A _2973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5755_ _1679_ _1678_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8543_ net235 net233 net199 _3994_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__and4b_1
X_4706_ net224 allocation.game.cactusMove.x_dist\[5\] vssd1 vssd1 vccd1 vccd1 _0633_
+ sky130_fd_sc_hd__or2_1
X_5686_ _1609_ _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__nand2b_1
X_8474_ net37 net43 _3356_ _3277_ vssd1 vssd1 vccd1 vccd1 _3927_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_20_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4637_ _0560_ _0566_ _0559_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7425_ net249 net252 vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__nand2_1
X_9516__301 vssd1 vssd1 vccd1 vccd1 _9516__301/HI net301 sky130_fd_sc_hd__conb_1
XFILLER_0_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4568_ net269 allocation.game.controller.v\[4\] _0505_ vssd1 vssd1 vccd1 vccd1 _0506_
+ sky130_fd_sc_hd__a21o_1
X_7356_ allocation.game.lcdOutput.tft.remainingDelayTicks\[19\] _2995_ vssd1 vssd1
+ vccd1 vccd1 _2996_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7287_ allocation.game.controller.init_module.delay_counter\[10\] _2946_ vssd1 vssd1
+ vccd1 vccd1 _2947_ sky130_fd_sc_hd__and2_1
X_4499_ allocation.game.scoreCounter.bcd_tens\[5\] vssd1 vssd1 vccd1 vccd1 _0439_
+ sky130_fd_sc_hd__inv_2
X_6307_ _1228_ _2131_ _2160_ _2162_ _2231_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__o2111ai_1
X_9026_ clknet_leaf_5_clk _0151_ net182 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6238_ _1328_ _1330_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__nor2_1
X_6169_ _2085_ _2093_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8078__A _0541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__6061__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5540_ _1439_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5471_ _1395_ _1394_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__and2b_1
X_7210_ allocation.game.dinoJump.count\[10\] allocation.game.dinoJump.count\[11\]
+ _2886_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8190_ _0652_ _0662_ _0651_ vssd1 vssd1 vccd1 vccd1 _3681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7141_ _2839_ _2843_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7072_ allocation.game.controller.drawBlock.x_start\[1\] _2772_ _2777_ allocation.game.controller.drawBlock.x_end\[1\]
+ _2790_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__a221o_1
X_6023_ _0723_ net102 _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4963__B _0708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout170_A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7974_ net278 net275 vssd1 vssd1 vccd1 vccd1 _3486_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout268_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6925_ _2690_ _2691_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7619__X _3181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout47 _3248_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_4
Xfanout36 _3263_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_2
X_6856_ _2642_ _2643_ _2644_ _2645_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__or4_2
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5807_ net87 _0905_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__and2_1
Xfanout58 _3218_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout69 _3208_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_4
X_6787_ allocation.game.cactus2size.clock_div_inst1.counter\[5\] allocation.game.cactus2size.clock_div_inst1.counter\[4\]
+ _2596_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5738_ _1660_ _1662_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__nand2_1
X_8526_ net56 _3298_ _3864_ net66 vssd1 vssd1 vccd1 vccd1 _3978_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8457_ _3345_ _3880_ vssd1 vssd1 vccd1 vccd1 _3910_ sky130_fd_sc_hd__nand2_1
X_5669_ _1591_ _1592_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__xnor2_1
X_8388_ _3476_ _3846_ _3842_ vssd1 vssd1 vccd1 vccd1 _3847_ sky130_fd_sc_hd__a21oi_1
X_7408_ _0420_ _3018_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__nand2_1
X_7339_ allocation.game.cactusHeight1\[2\] _2975_ _2982_ vssd1 vssd1 vccd1 vccd1 _0198_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9009_ net255 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__inv_2
XANTENNA__5985__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5942__B1 _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_X clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload17 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9292__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4971_ net78 _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nor2_4
X_6710_ allocation.game.cactus1size.clock_div_inst1.counter\[7\] allocation.game.cactus1size.clock_div_inst1.counter\[8\]
+ _2544_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__and3_1
X_7690_ allocation.game.lcdOutput.framebufferIndex\[5\] net47 vssd1 vssd1 vccd1 vccd1
+ _3252_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6641_ _2502_ _2503_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[24\]
+ sky130_fd_sc_hd__nor2_1
X_9360_ clknet_leaf_12_clk _0009_ net204 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_8311_ _3773_ _3775_ _3776_ vssd1 vssd1 vccd1 vccd1 _3777_ sky130_fd_sc_hd__or3b_1
X_6572_ allocation.game.cactusMove.count\[29\] allocation.game.cactusMove.count\[28\]
+ allocation.game.cactusMove.count\[31\] allocation.game.cactusMove.count\[30\] vssd1
+ vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5523_ _0918_ _1447_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__nand2_1
X_9291_ clknet_leaf_0_clk _0093_ net166 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8478__A2 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5454_ _0754_ _0821_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__xnor2_1
X_8242_ _2990_ _3720_ _3000_ vssd1 vssd1 vccd1 vccd1 _3721_ sky130_fd_sc_hd__a21o_1
X_8173_ net113 _2520_ _3609_ net101 _3598_ vssd1 vssd1 vccd1 vccd1 _3666_ sky130_fd_sc_hd__o221a_1
X_5385_ _1303_ _1305_ _1309_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__o21a_1
Xfanout204 net205 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
XANTENNA__5135__A _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7124_ _2830_ _2831_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_2
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_4
Xfanout226 allocation.game.cactusMove.pixel\[4\] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7055_ _2773_ _2774_ net236 vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__o21a_1
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
Xfanout248 allocation.game.lcdOutput.tft.initSeqCounter\[3\] vssd1 vssd1 vccd1 vccd1
+ net248 sky130_fd_sc_hd__buf_2
X_6006_ _1886_ _1887_ _1889_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7610__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7957_ _0496_ _0523_ vssd1 vssd1 vccd1 vccd1 _3470_ sky130_fd_sc_hd__or2_1
XANTENNA__5563__A_N net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7888_ allocation.game.controller.drawBlock.counter\[6\] _3420_ net94 vssd1 vssd1
+ vccd1 vccd1 _3424_ sky130_fd_sc_hd__o21ai_1
X_6908_ _2679_ _2680_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6839_ allocation.game.cactus2size.clock_div_inst0.counter\[9\] _2633_ vssd1 vssd1
+ vccd1 vccd1 _2634_ sky130_fd_sc_hd__and2_1
XANTENNA__7913__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9165__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9489_ clknet_leaf_3_clk _0389_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.r_idle
+ sky130_fd_sc_hd__dfxtp_1
X_8509_ _3337_ _3864_ net56 _3318_ vssd1 vssd1 vccd1 vccd1 _3961_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout86_X net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5455__A2 _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9423__Q allocation.game.controller.drawBlock.y_start\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5170_ _1074_ _1091_ _1093_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__or3b_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 gpio_in[2] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
XANTENNA__9038__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8860_ net38 _4304_ vssd1 vssd1 vccd1 vccd1 _4310_ sky130_fd_sc_hd__nor2_1
X_7811_ _3309_ _3369_ _3372_ net118 vssd1 vssd1 vccd1 vccd1 _3373_ sky130_fd_sc_hd__a211o_1
X_8791_ _4214_ _4216_ _4219_ net36 _4240_ vssd1 vssd1 vccd1 vccd1 _4241_ sky130_fd_sc_hd__a221o_1
X_4954_ _0877_ _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__and2_1
X_7742_ net66 net58 _3302_ vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9412_ clknet_leaf_13_clk _0321_ net210 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.wr
+ sky130_fd_sc_hd__dfstp_1
X_4885_ _0740_ _0742_ _0764_ _0781_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_28_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7673_ _3226_ _3234_ vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_41_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6624_ allocation.game.cactusMove.count\[18\] _2490_ net149 vssd1 vssd1 vccd1 vccd1
+ _2493_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9343_ clknet_leaf_2_clk _0275_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.game.score\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_6555_ net397 _2443_ _2445_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[17\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9274_ clknet_leaf_4_clk _0262_ net187 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.lfsr1\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_5506_ _0820_ _0822_ _0725_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__mux2_1
X_6486_ allocation.game.scoreCounter.clock_div.counter\[7\] _2391_ _2392_ _2400_ vssd1
+ vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__or4b_1
XANTENNA__8320__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8225_ allocation.game.lcdOutput.tft.remainingDelayTicks\[4\] _2985_ net454 vssd1
+ vssd1 vccd1 vccd1 _3710_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5437_ _1360_ _1361_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__nor2_1
X_8156_ net218 _3644_ vssd1 vssd1 vccd1 vccd1 _3654_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_39_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5368_ _1031_ _1292_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7107_ allocation.game.controller.init_module.delay_counter\[15\] allocation.game.controller.init_module.delay_counter\[14\]
+ allocation.game.controller.init_module.delay_counter\[13\] allocation.game.controller.init_module.delay_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__or4_1
X_8087_ net257 net77 _0627_ net206 vssd1 vssd1 vccd1 vccd1 _3592_ sky130_fd_sc_hd__o211a_1
XANTENNA__4908__S _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5299_ _1222_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8623__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7038_ _0425_ allocation.game.controller.init_module.idx\[2\] _2758_ vssd1 vssd1
+ vccd1 vccd1 _2759_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_48_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8989_ _4437_ vssd1 vssd1 vccd1 vccd1 _4438_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout46_A _3256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7239__B _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7898__B1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5125__A1 _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8075__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8086__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8814__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9330__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9480__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4670_ _0584_ _0599_ _0583_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9499__284 vssd1 vssd1 vccd1 vccd1 _9499__284/HI net284 sky130_fd_sc_hd__conb_1
XFILLER_0_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6340_ allocation.game.collision.dinoY\[0\] allocation.game.cactusHeight2\[0\] _2260_
+ net279 vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7165__A _0401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6271_ _2080_ _2096_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__nand2_1
X_5222_ _1141_ _1145_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__xnor2_2
X_8010_ net270 _3509_ vssd1 vssd1 vccd1 vccd1 _3520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5153_ _0805_ _0810_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__xnor2_1
X_5084_ _0893_ net64 _1008_ _0798_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__a22o_1
X_8912_ _4354_ _4361_ net44 vssd1 vssd1 vccd1 vccd1 _4362_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8843_ _4228_ _4248_ _4292_ _4227_ vssd1 vssd1 vccd1 vccd1 _4293_ sky130_fd_sc_hd__o211a_1
XANTENNA__4971__B _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5986_ net110 _0905_ _1865_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__a21o_1
X_8774_ _4212_ _4223_ net128 vssd1 vssd1 vccd1 vccd1 _4224_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _0798_ _0860_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__and2_1
X_7725_ _4454_ net126 _3286_ _3281_ vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4868_ _0771_ _0779_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__or2_1
X_7656_ _3212_ _3214_ _3216_ vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6607_ allocation.game.cactusMove.count\[12\] _2480_ vssd1 vssd1 vccd1 vccd1 _2482_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9326_ clknet_leaf_6_clk _0109_ net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_4799_ _0709_ net110 vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_31_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7587_ allocation.game.cactus2size.lfsr1\[1\] allocation.game.cactus2size.lfsr1\[0\]
+ allocation.game.cactus2size.clock_div_inst0.clk1 vssd1 vssd1 vccd1 vccd1 _3166_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6538_ net387 _2432_ _2434_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[11\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6469_ net232 _0446_ net234 vssd1 vssd1 vccd1 vccd1 _2386_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9257_ clknet_leaf_0_clk _0065_ net177 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8208_ _3689_ _3691_ _3697_ net207 net383 vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__o32a_1
X_9188_ clknet_leaf_15_clk _0250_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8139_ _0679_ _3626_ _3637_ net243 vssd1 vssd1 vccd1 vccd1 _3638_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9353__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7099__A1 allocation.game.controller.drawBlock.y_end\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7032__A_N allocation.game.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5840_ _1752_ _1753_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5771_ _0897_ _1695_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4722_ net112 _0648_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__nor2_1
X_8490_ _3918_ _3942_ _3940_ _3862_ vssd1 vssd1 vccd1 vccd1 _3943_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7510_ _0430_ net250 _3048_ _3054_ _3084_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__o32a_1
X_7441_ _0429_ net245 vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__nor2_1
XANTENNA__7607__B _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4653_ allocation.game.controller.drawBlock.y_start\[4\] allocation.game.controller.drawBlock.y_end\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9226__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4584_ net276 _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nand2_1
XANTENNA__7326__C net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7372_ _2998_ _3006_ net55 vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__a21oi_1
X_9111_ clknet_leaf_7_clk allocation.game.cactusMove.n_count\[5\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[5\] sky130_fd_sc_hd__dfrtp_1
X_6323_ _2244_ _2245_ _2246_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__and3_1
XANTENNA__8719__A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9042_ clknet_leaf_7_clk _0167_ net184 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_6254_ allocation.game.controller.drawBlock.counter\[15\] _2177_ vssd1 vssd1 vccd1
+ vccd1 _2179_ sky130_fd_sc_hd__nor2_1
XANTENNA__9376__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5205_ net83 _1126_ _1128_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6185_ _2108_ _2109_ _1943_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__a21boi_1
X_5136_ _1051_ _1055_ _1060_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__o21a_1
X_5067_ _0990_ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__nand2_2
X_8826_ _4217_ _4241_ _4275_ vssd1 vssd1 vccd1 vccd1 _4276_ sky130_fd_sc_hd__a21bo_1
X_5969_ _1847_ _1892_ _1891_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__o21ai_1
X_8757_ net34 _3284_ _4121_ _4207_ _4077_ vssd1 vssd1 vccd1 vccd1 _4208_ sky130_fd_sc_hd__o311a_1
X_7708_ _3269_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8688_ net52 _3603_ _4138_ vssd1 vssd1 vccd1 vccd1 _4139_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7639_ allocation.game.lcdOutput.framebufferIndex\[10\] net74 vssd1 vssd1 vccd1 vccd1
+ _3201_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9309_ clknet_leaf_3_clk _0269_ net191 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.lfsr1\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__8348__B net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8364__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8753__A1 _3219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9249__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9399__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8269__A0 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 allocation.game.cactus1size.clock_div_inst1.counter\[3\] vssd1 vssd1 vccd1
+ vccd1 net432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5898__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7990_ net81 net77 vssd1 vssd1 vccd1 vccd1 _3502_ sky130_fd_sc_hd__nand2_2
X_6941_ allocation.game.scoreCounter.clock_div.counter\[3\] _2396_ vssd1 vssd1 vccd1
+ vccd1 _2700_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6872_ allocation.game.cactusDist.clock_div_inst1.counter\[6\] _2655_ vssd1 vssd1
+ vccd1 vccd1 _2656_ sky130_fd_sc_hd__and2_1
X_8611_ _0614_ _2375_ net75 vssd1 vssd1 vccd1 vccd1 _4062_ sky130_fd_sc_hd__or3_1
X_5823_ _1730_ _1731_ _1747_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8542_ _3956_ _3985_ _3989_ _3993_ vssd1 vssd1 vccd1 vccd1 _3994_ sky130_fd_sc_hd__or4b_1
XFILLER_0_45_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5754_ _0990_ _1668_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4705_ net224 allocation.game.cactusMove.x_dist\[5\] vssd1 vssd1 vccd1 vccd1 _0632_
+ sky130_fd_sc_hd__nand2_1
X_5685_ _1565_ _1567_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__xnor2_1
X_8473_ _3908_ _3911_ _3923_ _3925_ _3271_ vssd1 vssd1 vccd1 vccd1 _3926_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout213_A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4636_ _0564_ _0565_ _0562_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7424_ net251 allocation.game.lcdOutput.tft.initSeqCounter\[1\] vssd1 vssd1 vccd1
+ vccd1 _3041_ sky130_fd_sc_hd__nand2_1
X_7355_ allocation.game.lcdOutput.tft.remainingDelayTicks\[18\] _2994_ vssd1 vssd1
+ vccd1 vccd1 _2995_ sky130_fd_sc_hd__or2_1
X_4567_ _0487_ _0502_ _0504_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__a21oi_1
X_6306_ _1328_ _2129_ _2163_ _2128_ _2230_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__o221a_1
X_7286_ _2927_ _2945_ _2946_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__nor3_1
X_4498_ allocation.game.scoreCounter.clock_div.slow_clk vssd1 vssd1 vccd1 vccd1 _0438_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9025_ clknet_leaf_5_clk _0150_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6237_ _2130_ _2161_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__or2_1
XANTENNA__4983__Y _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6168_ _2082_ _2084_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__or2_1
X_5119_ _1009_ _1043_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__or2_1
X_6099_ _2020_ _2021_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8735__B2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8735__A1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8809_ _4257_ _4258_ vssd1 vssd1 vccd1 vccd1 _4259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5511__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9071__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9426__Q allocation.game.controller.drawBlock.y_start\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5470_ _0864_ _1391_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7140_ allocation.game.lcdOutput.framebufferIndex\[15\] net125 allocation.game.lcdOutput.framebufferIndex\[12\]
+ allocation.game.lcdOutput.framebufferIndex\[13\] vssd1 vssd1 vccd1 vccd1 _2843_
+ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_18_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7071_ allocation.game.controller.drawBlock.y_end\[1\] _2779_ _2787_ allocation.game.controller.drawBlock.y_start\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__a22o_1
XANTENNA__9161__Q allocation.game.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6022_ _0716_ _0907_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__nand2_1
XANTENNA__9414__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5421__A _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7973_ _3480_ _3481_ _3485_ net197 net409 vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__o32a_1
X_6924_ net404 _2689_ net155 vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_1_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout37 _3261_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_4
X_6855_ allocation.game.cactusDist.clock_div_inst1.counter\[11\] allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ allocation.game.cactusDist.clock_div_inst1.counter\[13\] allocation.game.cactusDist.clock_div_inst1.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__or4_1
X_5806_ _1678_ _1679_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__xnor2_1
Xfanout48 _3236_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
X_6786_ allocation.game.cactus2size.clock_div_inst1.counter\[4\] _2596_ allocation.game.cactus2size.clock_div_inst1.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__a21oi_1
Xfanout59 _3218_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5737_ net63 _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__nand2_1
X_8525_ net126 _3311_ _3971_ _3976_ _3271_ vssd1 vssd1 vccd1 vccd1 _3977_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8456_ net43 net34 _3356_ _3277_ vssd1 vssd1 vccd1 vccd1 _3909_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7407_ _3027_ _3028_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__and2_1
X_5668_ _1592_ _1591_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__and2b_1
X_8387_ allocation.game.controller.v\[1\] allocation.game.controller.v\[0\] allocation.game.controller.v\[2\]
+ vssd1 vssd1 vccd1 vccd1 _3846_ sky130_fd_sc_hd__o21ai_1
X_4619_ _0547_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__nand2b_1
X_5599_ _1471_ _1522_ _1523_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7338_ _2978_ _2981_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7269_ net470 _2933_ net122 vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9008_ allocation.game.controller.state\[6\] vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__9094__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5331__A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8642__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5942__A1 _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5942__B2 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6498__A2 allocation.game.dinoJump.dinoMovement vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9437__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6337__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4970_ _0591_ _0697_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__nand2_4
XANTENNA__8552__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6640_ allocation.game.cactusMove.count\[24\] _2501_ net150 vssd1 vssd1 vccd1 vccd1
+ _2503_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6571_ allocation.game.cactusMove.count\[25\] allocation.game.cactusMove.count\[24\]
+ allocation.game.cactusMove.count\[27\] allocation.game.cactusMove.count\[26\] vssd1
+ vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__or4_1
X_8310_ _2280_ net100 _2411_ net274 net198 vssd1 vssd1 vccd1 vccd1 _3776_ sky130_fd_sc_hd__o221a_1
X_5522_ _1445_ _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9290_ clknet_leaf_0_clk _0092_ net166 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8241_ allocation.game.lcdOutput.tft.remainingDelayTicks\[10\] _2989_ allocation.game.lcdOutput.tft.remainingDelayTicks\[11\]
+ vssd1 vssd1 vccd1 vccd1 _3720_ sky130_fd_sc_hd__o21ai_1
X_5453_ _1325_ _1375_ _1376_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__and3_1
X_8172_ _3597_ _3663_ _3665_ net203 net451 vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__o32a_1
X_5384_ _1307_ _1308_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nor2_1
Xfanout205 net216 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
XANTENNA__8635__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7123_ allocation.game.lcdOutput.framebufferIndex\[4\] net127 _0453_ allocation.game.lcdOutput.framebufferIndex\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout238 allocation.game.controller.block_done vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout216 allocation.game.cactus1size.clock_div_inst0.reset vssd1 vssd1 vccd1 vccd1
+ net216 sky130_fd_sc_hd__buf_2
Xfanout227 allocation.game.cactusMove.pixel\[3\] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7054_ allocation.game.controller.drawBlock.idx\[3\] allocation.game.controller.drawBlock.idx\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__nand2b_1
Xfanout249 allocation.game.lcdOutput.tft.initSeqCounter\[3\] vssd1 vssd1 vccd1 vccd1
+ net249 sky130_fd_sc_hd__buf_2
XANTENNA_fanout280_A allocation.game.collision.dinoY\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_6005_ _1907_ _1927_ _1928_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__nand3_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7956_ allocation.game.controller.drawBlock.y_start\[0\] net204 _3468_ _3469_ vssd1
+ vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7887_ allocation.game.controller.drawBlock.counter\[6\] _3420_ vssd1 vssd1 vccd1
+ vccd1 _3423_ sky130_fd_sc_hd__and2_1
X_6907_ allocation.game.cactusDist.clock_div_inst0.counter\[3\] _2678_ net155 vssd1
+ vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6838_ net160 _2632_ _2633_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__nor3_1
XFILLER_0_18_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8508_ _3282_ _3341_ _3959_ _3958_ vssd1 vssd1 vccd1 vccd1 _3960_ sky130_fd_sc_hd__a31o_1
X_6769_ allocation.game.cactus2size.clock_div_inst1.counter\[0\] _2586_ allocation.game.cactus2size.clock_div_inst1.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9488_ clknet_leaf_11_clk allocation.game.cactusMove.n_pixel\[8\] net201 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.pixel\[8\] sky130_fd_sc_hd__dfstp_1
X_8439_ _3318_ _3864_ vssd1 vssd1 vccd1 vccd1 _3892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6157__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9529__323 vssd1 vssd1 vccd1 vccd1 net323 _9529__323/LO sky130_fd_sc_hd__conb_1
XFILLER_0_38_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7716__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9501__286 vssd1 vssd1 vccd1 vccd1 _9501__286/HI net286 sky130_fd_sc_hd__conb_1
XFILLER_0_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6340__A1 allocation.game.collision.dinoY\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7451__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 nrst vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_2
X_7810_ _3305_ _3369_ _3371_ vssd1 vssd1 vccd1 vccd1 _3372_ sky130_fd_sc_hd__a21oi_1
X_8790_ net36 _4219_ _4238_ _4239_ _4221_ vssd1 vssd1 vccd1 vccd1 _4240_ sky130_fd_sc_hd__o221a_1
X_4953_ _0870_ _0876_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__nand2_1
X_7741_ net66 net58 vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__nand2_1
X_7672_ _3223_ net50 _3225_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9411_ clknet_leaf_13_clk _0398_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.init_done
+ sky130_fd_sc_hd__dfrtp_1
X_4884_ _0760_ _0808_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__xnor2_4
X_6623_ allocation.game.cactusMove.count\[18\] _2490_ vssd1 vssd1 vccd1 vccd1 _2492_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_41_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9342_ clknet_leaf_1_clk _0274_ net165 vssd1 vssd1 vccd1 vccd1 allocation.game.game.score\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_6554_ allocation.game.dinoJump.dinoDelay\[17\] _2443_ net90 vssd1 vssd1 vccd1 vccd1
+ _2445_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout126_A allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6485_ allocation.game.scoreCounter.clock_div.counter\[16\] allocation.game.scoreCounter.clock_div.counter\[15\]
+ allocation.game.scoreCounter.clock_div.counter\[0\] vssd1 vssd1 vccd1 vccd1 _2400_
+ sky130_fd_sc_hd__and3_1
X_5505_ _0806_ _1429_ _0813_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__mux2_1
X_9273_ clknet_leaf_2_clk _0052_ net181 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5874__A2_N net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8224_ _3033_ _3708_ _3709_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5436_ _1353_ _1356_ _1359_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_39_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8155_ _0415_ _0618_ net218 vssd1 vssd1 vccd1 vccd1 _3653_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_39_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5367_ _1290_ _1291_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7106_ allocation.game.controller.init_module.delay_counter\[9\] _2817_ allocation.game.controller.init_module.delay_counter\[11\]
+ allocation.game.controller.init_module.delay_counter\[10\] vssd1 vssd1 vccd1 vccd1
+ _2818_ sky130_fd_sc_hd__o211a_1
X_8086_ net257 _0682_ vssd1 vssd1 vccd1 vccd1 _3591_ sky130_fd_sc_hd__nand2_1
X_5298_ _1216_ _1220_ _1221_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__nand3_1
X_7037_ net4 _2757_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_21_clk_X clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9132__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8988_ net46 _4149_ _4169_ _4431_ vssd1 vssd1 vccd1 vccd1 _4437_ sky130_fd_sc_hd__or4_1
X_7939_ _0424_ _0399_ _3458_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9282__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6322__A1 _4459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8075__A1 _0541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6270_ _2098_ _2194_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__or2_1
X_5221_ _1145_ _1141_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5152_ _0806_ _0810_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9155__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5083_ _0924_ net60 vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__xor2_1
X_8911_ _4298_ _4299_ _4358_ _4360_ _4356_ vssd1 vssd1 vccd1 vccd1 _4361_ sky130_fd_sc_hd__o32a_1
XFILLER_0_21_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8842_ _4282_ _4287_ _4288_ _4291_ vssd1 vssd1 vccd1 vccd1 _4292_ sky130_fd_sc_hd__and4b_1
X_8773_ _4458_ _3486_ vssd1 vssd1 vccd1 vccd1 _4223_ sky130_fd_sc_hd__or2_1
X_5985_ net103 _0904_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__nor2_1
X_7724_ _2861_ _3285_ vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout243_A allocation.game.controller.state\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4936_ _0798_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4867_ _0783_ _0784_ _0786_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__o21ai_2
X_7655_ _3214_ _3216_ vssd1 vssd1 vccd1 vccd1 _3217_ sky130_fd_sc_hd__nand2_1
X_6606_ _2480_ _2481_ _2462_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[11\]
+ sky130_fd_sc_hd__and3b_1
X_7586_ allocation.game.cactus2size.lfsr1\[0\] _3164_ _3165_ vssd1 vssd1 vccd1 vccd1
+ _0262_ sky130_fd_sc_hd__o21ai_1
X_9325_ clknet_leaf_6_clk _0108_ net174 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_4798_ _0720_ _0721_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_31_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6537_ allocation.game.dinoJump.dinoDelay\[11\] _2432_ net90 vssd1 vssd1 vccd1 vccd1
+ _2434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6468_ _2372_ _2384_ vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__nor2_1
X_9256_ clknet_leaf_0_clk _0064_ net176 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8207_ net101 _3695_ _3696_ net113 net205 vssd1 vssd1 vccd1 vccd1 _3697_ sky130_fd_sc_hd__o221ai_2
X_9187_ clknet_leaf_15_clk _0249_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataDc
+ sky130_fd_sc_hd__dfxtp_1
X_6399_ allocation.game.game.score\[2\] _2321_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7803__B net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5419_ _0938_ _1201_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__nand2_1
X_8138_ net105 _3626_ vssd1 vssd1 vccd1 vccd1 _3637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8069_ net263 _2412_ _3576_ net244 _3501_ vssd1 vssd1 vccd1 vccd1 _3577_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_6_Left_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9028__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4609__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5770_ _1692_ _1693_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__xnor2_1
X_9507__292 vssd1 vssd1 vccd1 vccd1 _9507__292/HI net292 sky130_fd_sc_hd__conb_1
X_4721_ net121 _0647_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nand2_1
X_4652_ _0580_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__nand2b_1
XANTENNA__7176__A _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7440_ _3056_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__inv_2
X_9110_ clknet_leaf_7_clk allocation.game.cactusMove.n_count\[4\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[4\] sky130_fd_sc_hd__dfrtp_1
X_4583_ _0472_ _0479_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__nor2_1
X_7371_ net366 _2997_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__nand2_1
X_6322_ _4459_ _2240_ _2243_ net265 vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9041_ clknet_leaf_7_clk _0166_ net184 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_6253_ allocation.game.controller.drawBlock.counter\[15\] _2177_ vssd1 vssd1 vccd1
+ vccd1 _2178_ sky130_fd_sc_hd__and2_1
X_5204_ net82 _1126_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__nand3_1
XANTENNA__4848__A1 _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6184_ _1941_ _1942_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_48_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5135_ _1052_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout193_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5066_ net82 _0820_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__or2_1
X_8825_ _4272_ _4274_ _3931_ vssd1 vssd1 vccd1 vccd1 _4275_ sky130_fd_sc_hd__or3b_1
X_5968_ _1847_ _1891_ _1892_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__or3_1
X_8756_ _4147_ _4178_ _4206_ vssd1 vssd1 vccd1 vccd1 _4207_ sky130_fd_sc_hd__a21bo_1
X_4919_ _0837_ _0839_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4784__B1 _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7707_ net127 net35 _3268_ net39 vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__a31o_1
X_5899_ _0761_ _0907_ _1822_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__a21o_1
X_8687_ net59 _3607_ vssd1 vssd1 vccd1 vccd1 _4138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7638_ net74 vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7569_ _3155_ _3156_ allocation.game.lcdOutput.tft.spi.counter\[0\] vssd1 vssd1 vccd1
+ vccd1 _3157_ sky130_fd_sc_hd__mux2_1
XANTENNA__9320__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9308_ clknet_leaf_3_clk _0268_ net191 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.lfsr1\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9239_ clknet_leaf_22_clk _0023_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5053__B _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9470__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout61_X net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9402__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5898__B _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9003__X _4452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6940_ _2396_ net91 _2699_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__and3b_1
X_6871_ net159 _2654_ _2655_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__nor3_1
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8610_ net225 net69 vssd1 vssd1 vccd1 vccd1 _4061_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5822_ _1745_ _1746_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5753_ _0819_ _1669_ _1677_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__a21bo_1
X_8541_ _3953_ _3965_ _3975_ _3992_ vssd1 vssd1 vccd1 vccd1 _3993_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4704_ _0629_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__nand2_1
XANTENNA__5419__A _0938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9343__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5684_ _1605_ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__nor2_1
X_8472_ net45 _3357_ _3924_ _3274_ vssd1 vssd1 vccd1 vccd1 _3925_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_20_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4635_ allocation.game.controller.drawBlock.x_end\[1\] allocation.game.controller.drawBlock.x_start\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__xnor2_4
XANTENNA__5715__C1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7423_ net251 net252 vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__and2_1
X_4566_ net269 allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__xnor2_4
X_7354_ allocation.game.lcdOutput.tft.remainingDelayTicks\[17\] allocation.game.lcdOutput.tft.remainingDelayTicks\[16\]
+ _2993_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6305_ _2127_ _2164_ _2165_ _2124_ _2229_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__o221a_1
X_7285_ allocation.game.controller.init_module.delay_counter\[9\] allocation.game.controller.init_module.delay_counter\[8\]
+ _2942_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__and3_1
XANTENNA__5154__A _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4497_ allocation.game.cactusHeight2\[0\] vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9024_ allocation.game.lcdOutput.tft.frameBufferLowNibble vssd1 vssd1 vccd1 vccd1
+ _0149_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9493__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6236_ _1327_ _2129_ _1282_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__a21oi_1
X_6167_ _2089_ _2091_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__and2_1
X_5118_ _1014_ _1041_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__xnor2_1
X_6098_ _0741_ net124 vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__nor2_1
X_5049_ net73 _0754_ _0952_ _0954_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8808_ net40 _4256_ vssd1 vssd1 vccd1 vccd1 _4258_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8739_ _4181_ _4189_ vssd1 vssd1 vccd1 vccd1 _4190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8974__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9216__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9366__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7070_ allocation.game.controller.init_module.idx\[0\] allocation.game.controller.init_module.idx\[1\]
+ _0426_ _2758_ _2756_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__a41o_1
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6021_ _0715_ _0908_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7972_ net279 net139 _3484_ allocation.game.controller.state\[4\] vssd1 vssd1 vccd1
+ vccd1 _3485_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6923_ allocation.game.cactusDist.clock_div_inst0.counter\[9\] _2689_ vssd1 vssd1
+ vccd1 vccd1 _2690_ sky130_fd_sc_hd__and2_1
XANTENNA__9395__RESET_B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout38 _3260_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_2
XANTENNA__7925__B1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6854_ allocation.game.cactusDist.clock_div_inst1.counter\[7\] allocation.game.cactusDist.clock_div_inst1.counter\[6\]
+ allocation.game.cactusDist.clock_div_inst1.counter\[9\] allocation.game.cactusDist.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout156_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout49 _3236_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_2
X_5805_ _1729_ _1728_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__and2b_1
X_6785_ allocation.game.cactus2size.clock_div_inst1.counter\[4\] _2596_ _2598_ vssd1
+ vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__o21a_1
X_5736_ _1658_ _1659_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__xnor2_1
X_8524_ _3975_ _3973_ vssd1 vssd1 vccd1 vccd1 _3976_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8455_ _3326_ _3906_ _3907_ _3360_ vssd1 vssd1 vccd1 vccd1 _3908_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5667_ _1545_ _1546_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__xnor2_1
X_4618_ allocation.game.controller.drawBlock.x_end\[6\] allocation.game.controller.drawBlock.x_start\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7406_ _0420_ _3026_ vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__nand2_1
X_8386_ _3841_ _3845_ _3843_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__a21oi_1
X_5598_ _1461_ _1463_ _1470_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__nor3_1
X_4549_ net273 allocation.game.controller.v\[3\] vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__nand2_1
X_7337_ _2973_ _2977_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__nor2_1
X_7268_ allocation.game.controller.init_module.delay_counter\[3\] _2933_ vssd1 vssd1
+ vccd1 vccd1 _2935_ sky130_fd_sc_hd__and2_1
X_9007_ net241 vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__clkbuf_1
X_6219_ _1177_ _1232_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__xnor2_1
XANTENNA__9239__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7199_ net148 _2882_ _0472_ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout69_A _3208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9389__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9065__RESET_B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8642__B net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4898__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4681__A2 allocation.game.dinoJump.dinoMovement vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7168__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6570_ allocation.game.cactusMove.count\[19\] allocation.game.cactusMove.count\[18\]
+ allocation.game.cactusMove.count\[17\] allocation.game.cactusMove.count\[16\] vssd1
+ vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_27_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5521_ _0778_ _0888_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8240_ net54 _3719_ _3036_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5452_ _1325_ _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8171_ _3664_ vssd1 vssd1 vccd1 vccd1 _3665_ sky130_fd_sc_hd__inv_2
X_5383_ _1290_ _1306_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7122_ allocation.game.lcdOutput.framebufferIndex\[4\] allocation.game.lcdOutput.framebufferIndex\[5\]
+ net127 _0453_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__and4_1
Xfanout206 net207 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
X_7053_ allocation.game.controller.drawBlock.idx\[0\] _0444_ allocation.game.controller.drawBlock.idx\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__or3_1
Xfanout228 allocation.game.cactusMove.pixel\[3\] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_1
Xfanout217 allocation.game.cactusMove.pixel\[8\] vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
XANTENNA_clkload10_A clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6004_ _1907_ _1927_ _1928_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__and3_1
X_7955_ allocation.game.collision.dinoY\[0\] net163 _3464_ _3467_ vssd1 vssd1 vccd1
+ vccd1 _3469_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7886_ net94 _3421_ _3422_ net108 allocation.game.controller.drawBlock.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a32o_1
X_6906_ allocation.game.cactusDist.clock_div_inst0.counter\[3\] _2678_ vssd1 vssd1
+ vccd1 vccd1 _2679_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_46_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6837_ allocation.game.cactus2size.clock_div_inst0.counter\[7\] allocation.game.cactus2size.clock_div_inst0.counter\[8\]
+ _2629_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8507_ _0401_ net132 net130 _0442_ vssd1 vssd1 vccd1 vccd1 _3959_ sky130_fd_sc_hd__and4_1
X_6768_ allocation.game.cactus2size.clock_div_inst1.counter\[3\] allocation.game.cactus2size.clock_div_inst1.counter\[5\]
+ allocation.game.cactus2size.clock_div_inst1.counter\[4\] allocation.game.cactus2size.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__or4b_1
X_9487_ clknet_leaf_11_clk allocation.game.cactusMove.n_pixel\[7\] net201 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.pixel\[7\] sky130_fd_sc_hd__dfrtp_1
X_5719_ _0915_ _1643_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__nor2_1
X_6699_ allocation.game.cactus1size.clock_div_inst1.counter\[4\] _2539_ net158 vssd1
+ vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5607__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5688__A1 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8438_ _3888_ _3890_ vssd1 vssd1 vccd1 vccd1 _3891_ sky130_fd_sc_hd__nand2_1
X_8369_ _3580_ _3816_ _0541_ vssd1 vssd1 vccd1 vccd1 _3831_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9061__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9404__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9536__317 vssd1 vssd1 vccd1 vccd1 _9536__317/HI net317 sky130_fd_sc_hd__conb_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5332__A_N _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8563__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4952_ _0870_ _0876_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__or2_1
X_7740_ net99 net74 vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6800__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4883_ _0739_ _0763_ _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__a21oi_4
X_7671_ _3230_ _3232_ vssd1 vssd1 vccd1 vccd1 _3233_ sky130_fd_sc_hd__and2_1
X_6622_ _2490_ _2491_ _2462_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[17\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9410_ clknet_leaf_17_clk _0320_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_41_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9084__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6553_ _2443_ _2444_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[16\]
+ sky130_fd_sc_hd__nor2_1
X_9341_ clknet_leaf_1_clk _0273_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.game.score\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_6484_ allocation.game.scoreCounter.clock_div.counter\[6\] _2398_ vssd1 vssd1 vccd1
+ vccd1 _2399_ sky130_fd_sc_hd__and2_1
X_5504_ _0729_ _0795_ net71 _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__a31o_1
X_9272_ clknet_leaf_2_clk _0051_ net176 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_8223_ allocation.game.lcdOutput.tft.remainingDelayTicks\[4\] _2985_ vssd1 vssd1
+ vccd1 vccd1 _3709_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout119_A _3181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5435_ _1353_ _1356_ _1359_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8608__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8154_ _0618_ _2313_ vssd1 vssd1 vccd1 vccd1 _3652_ sky130_fd_sc_hd__nand2_1
X_5366_ _1283_ _1287_ _1289_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__or3_1
X_7105_ allocation.game.controller.init_module.delay_counter\[7\] allocation.game.controller.init_module.delay_counter\[6\]
+ allocation.game.controller.init_module.delay_counter\[8\] vssd1 vssd1 vccd1 vccd1
+ _2817_ sky130_fd_sc_hd__o21a_1
X_8085_ allocation.game.controller.drawBlock.x_end\[0\] net206 _3590_ vssd1 vssd1
+ vccd1 vccd1 _0336_ sky130_fd_sc_hd__o21a_1
X_5297_ _1216_ _1220_ _1221_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7036_ allocation.game.controller.init_module.idx\[3\] allocation.game.controller.init_module.idx\[5\]
+ allocation.game.controller.init_module.idx\[4\] vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_48_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8987_ _4425_ _4426_ _4428_ _4424_ _4435_ vssd1 vssd1 vccd1 vccd1 _4436_ sky130_fd_sc_hd__o221a_1
X_7938_ _0695_ _2826_ _0424_ vssd1 vssd1 vccd1 vccd1 _3458_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9427__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7869_ net94 net108 allocation.game.controller.drawBlock.counter\[0\] vssd1 vssd1
+ vccd1 vccd1 _0300_ sky130_fd_sc_hd__mux2_1
XANTENNA__8544__B1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8935__X _0392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7727__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5220_ _1143_ _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5151_ _1074_ _1075_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__or2_1
X_5082_ _1005_ _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8910_ _4322_ _4358_ _4359_ vssd1 vssd1 vccd1 vccd1 _4360_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8293__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8841_ net38 _4279_ _4284_ net44 _4286_ vssd1 vssd1 vccd1 vccd1 _4291_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8772_ net268 _4212_ vssd1 vssd1 vccd1 vccd1 _4222_ sky130_fd_sc_hd__xnor2_1
X_5984_ _0723_ net102 _1865_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__or3b_1
X_7723_ _3283_ _3284_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__or2_1
X_4935_ _0858_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__xnor2_1
X_4866_ _0732_ _0790_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7654_ _3205_ _3215_ vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__and2b_1
X_6605_ allocation.game.cactusMove.count\[9\] allocation.game.cactusMove.count\[10\]
+ _2475_ allocation.game.cactusMove.count\[11\] vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__a31o_1
X_4797_ _0720_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__nor2_2
X_7585_ allocation.game.cactus2size.lfsr1\[0\] _3164_ net144 vssd1 vssd1 vccd1 vccd1
+ _3165_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9324_ clknet_leaf_6_clk _0107_ net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6536_ _2432_ _2433_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[10\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6467_ _2342_ _2349_ _2356_ _2344_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__o31a_1
X_9255_ clknet_leaf_0_clk _0063_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_8206_ allocation.game.cactusMove.pixel\[7\] _0623_ vssd1 vssd1 vccd1 vccd1 _3696_
+ sky130_fd_sc_hd__xor2_1
X_9186_ clknet_leaf_15_clk net351 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataShift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_6398_ allocation.game.game.score\[1\] allocation.game.game.score\[0\] vssd1 vssd1
+ vccd1 vccd1 _2321_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_7_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5418_ _1341_ _1342_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__and2_1
X_8137_ _3627_ _3629_ _3636_ net207 net411 vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__o32a_1
X_5349_ _1270_ _1272_ _1273_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8068_ net139 _3573_ _3574_ _3575_ vssd1 vssd1 vccd1 vccd1 _3576_ sky130_fd_sc_hd__a31o_1
X_7019_ allocation.game.scoreCounter.bcd_tens\[6\] allocation.game.scoreCounter.bcd_tens\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8650__B net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9261__RESET_B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4609__A2 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9103__SET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8560__B _3609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4720_ net142 _0646_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4651_ allocation.game.controller.drawBlock.y_end\[5\] allocation.game.controller.drawBlock.y_start\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_25_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_clk_X clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4582_ _0501_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7370_ _2996_ _3005_ net54 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__a21oi_1
X_6321_ net259 net263 vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9040_ clknet_leaf_7_clk _0165_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__9122__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6252_ _2112_ _2113_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7623__C net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5203_ _1071_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6183_ _1982_ _2107_ _1981_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__o21bai_1
X_5134_ _1057_ _1058_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__and2b_1
XANTENNA__9272__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5065_ net83 _0820_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8747__B1 net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8824_ _3305_ _3919_ _4273_ _3874_ vssd1 vssd1 vccd1 vccd1 _4274_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8470__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5967_ _1843_ _1844_ _1846_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__o21ba_1
X_8755_ net111 _0675_ _4180_ _4205_ _0669_ vssd1 vssd1 vccd1 vccd1 _4206_ sky130_fd_sc_hd__o311a_1
X_4918_ _0797_ _0841_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5981__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7706_ _3252_ net42 vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__nor2_1
X_8686_ net59 _3607_ _4124_ _4136_ vssd1 vssd1 vccd1 vccd1 _4137_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _0762_ _0908_ _1822_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__or3b_1
X_7637_ allocation.game.lcdOutput.framebufferIndex\[10\] _3187_ _3193_ _3198_ vssd1
+ vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__a31o_1
X_4849_ _0760_ net88 _0771_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__mux2_2
X_7568_ allocation.game.lcdOutput.tft.spi.dataShift\[4\] allocation.game.lcdOutput.tft.spi.dataShift\[5\]
+ allocation.game.lcdOutput.tft.spi.dataShift\[6\] allocation.game.lcdOutput.tft.spi.dataShift\[7\]
+ allocation.game.lcdOutput.tft.spi.counter\[2\] allocation.game.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__mux4_1
X_9307_ clknet_leaf_21_clk _0080_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_6519_ _2421_ _2422_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[4\]
+ sky130_fd_sc_hd__nor2_1
X_7499_ _3075_ _3083_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9238_ clknet_leaf_22_clk _0022_ net178 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout99_A _3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9169_ clknet_leaf_15_clk _0231_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8380__B _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9295__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7740__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8977__B1 _3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6870_ allocation.game.cactusDist.clock_div_inst1.counter\[5\] allocation.game.cactusDist.clock_div_inst1.counter\[4\]
+ _2651_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__and3_1
XANTENNA__8571__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5821_ _1730_ _1731_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_33_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5752_ _1676_ _1675_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__nand2b_1
X_8540_ _3270_ _3883_ _3991_ _3990_ vssd1 vssd1 vccd1 vccd1 _3992_ sky130_fd_sc_hd__o31a_1
XANTENNA__5963__B1 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4703_ net222 allocation.game.cactusMove.x_dist\[6\] vssd1 vssd1 vccd1 vccd1 _0630_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5683_ _1606_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__and2b_1
X_8471_ net35 _3361_ vssd1 vssd1 vccd1 vccd1 _3924_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4634_ allocation.game.controller.drawBlock.x_end\[0\] allocation.game.controller.drawBlock.x_start\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7422_ _3020_ _3031_ _3037_ _3039_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__a31o_2
XANTENNA__4610__Y _0541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4565_ allocation.game.controller.v\[4\] net270 vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__nand2b_1
X_7353_ allocation.game.lcdOutput.tft.remainingDelayTicks\[15\] _2992_ vssd1 vssd1
+ vccd1 vccd1 _2993_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6304_ allocation.game.controller.drawBlock.counter\[20\] _2168_ _2228_ _2166_ _2167_
+ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__o2111a_1
X_7284_ allocation.game.controller.init_module.delay_counter\[8\] _2942_ allocation.game.controller.init_module.delay_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__a21oi_1
X_4496_ allocation.game.cactusHeight1\[0\] vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9023_ net254 vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__inv_2
X_6235_ _1228_ _1230_ _1280_ _2130_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4993__B net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6166_ _2082_ _2090_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__nor2_1
X_5117_ _1041_ _1014_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__and2b_1
X_6097_ _1946_ _2019_ _2021_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__and3_1
X_5048_ _0964_ _0966_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__nand2b_1
X_9523__308 vssd1 vssd1 vccd1 vccd1 _9523__308/HI net308 sky130_fd_sc_hd__conb_1
X_8807_ net40 _4256_ vssd1 vssd1 vccd1 vccd1 _4257_ sky130_fd_sc_hd__nor2_1
X_6999_ allocation.game.bcd_ones\[2\] allocation.game.bcd_ones\[1\] vssd1 vssd1 vccd1
+ vccd1 _2736_ sky130_fd_sc_hd__and2b_1
X_8738_ net111 _4180_ vssd1 vssd1 vccd1 vccd1 _4189_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8669_ net131 _3312_ _3356_ net128 vssd1 vssd1 vccd1 vccd1 _4120_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5511__C _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8566__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6020_ _0769_ _0894_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_3_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__8285__B net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7971_ net140 _3482_ vssd1 vssd1 vccd1 vccd1 _3484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6922_ net161 _2688_ _2689_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9310__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6853_ allocation.game.cactusDist.clock_div_inst1.counter\[3\] allocation.game.cactusDist.clock_div_inst1.counter\[5\]
+ allocation.game.cactusDist.clock_div_inst1.counter\[4\] allocation.game.cactusDist.clock_div_inst1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__or4b_1
X_5804_ _1675_ _1676_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout39 _3260_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_2
X_6784_ allocation.game.cactus2size.clock_div_inst1.counter\[4\] _2596_ net162 vssd1
+ vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9460__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5735_ _1658_ _1659_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__nand2b_1
X_8523_ _3880_ _3961_ _3974_ vssd1 vssd1 vccd1 vccd1 _3975_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5666_ _1121_ _1579_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__o21ai_1
X_8454_ net118 _3289_ _3321_ _3893_ vssd1 vssd1 vccd1 vccd1 _3907_ sky130_fd_sc_hd__or4_1
XANTENNA__8350__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4617_ allocation.game.controller.drawBlock.x_start\[6\] allocation.game.controller.drawBlock.x_end\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7405_ allocation.game.lcdOutput.tft.state\[0\] _3025_ vssd1 vssd1 vccd1 vccd1 _3027_
+ sky130_fd_sc_hd__nand2_1
X_8385_ _3840_ _3844_ vssd1 vssd1 vccd1 vccd1 _3845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5597_ _1519_ _1521_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__nor2_1
X_4548_ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__or2_2
X_7336_ allocation.game.cactusHeight1\[1\] _2976_ _2979_ vssd1 vssd1 vccd1 vccd1 _0197_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout104_X net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7267_ _2933_ _2934_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__nor2_1
X_4479_ net243 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6218_ _2140_ _2142_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__xnor2_1
X_9006_ net282 _4452_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__nor2_1
X_7198_ _2878_ _2880_ _2881_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__and3_1
X_6149_ _2070_ _2073_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__nand2_1
XANTENNA__7613__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7916__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9034__RESET_B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8341__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7852__A0 allocation.game.controller.block_done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9333__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9010__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9483__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5520_ net71 _0885_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5451_ net61 _1324_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__or2_1
X_8170_ net81 net77 _0657_ vssd1 vssd1 vccd1 vccd1 _3664_ sky130_fd_sc_hd__mux2_1
X_5382_ _1290_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7121_ allocation.game.lcdOutput.framebufferIndex\[4\] _2828_ vssd1 vssd1 vccd1 vccd1
+ _0409_ sky130_fd_sc_hd__xnor2_1
Xfanout207 net216 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
X_7052_ _2770_ _2771_ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__nor2_2
Xfanout229 allocation.game.cactusMove.pixel\[2\] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
Xfanout218 allocation.game.cactusMove.pixel\[8\] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6003_ _1883_ _1926_ _1925_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__a21o_1
XANTENNA__7071__B2 allocation.game.controller.drawBlock.y_start\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7071__A1 allocation.game.controller.drawBlock.y_end\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_7954_ allocation.game.controller.state\[4\] net242 _3463_ vssd1 vssd1 vccd1 vccd1
+ _3468_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout266_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6905_ net161 _2677_ _2678_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__nor3_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7885_ allocation.game.controller.drawBlock.counter\[4\] _3415_ allocation.game.controller.drawBlock.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3422_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_18_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6836_ allocation.game.cactus2size.clock_div_inst0.counter\[7\] _2629_ allocation.game.cactus2size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__a21oi_1
X_6767_ net334 _2583_ _2585_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__a21oi_1
XANTENNA__7646__Y _3208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5718_ _0906_ _0913_ _1642_ net124 net78 vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8506_ net37 net42 _3957_ _3277_ vssd1 vssd1 vccd1 vccd1 _3958_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9486_ clknet_leaf_10_clk allocation.game.cactusMove.n_pixel\[6\] net196 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.pixel\[6\] sky130_fd_sc_hd__dfstp_1
X_6698_ _0447_ _2537_ _2540_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__a21oi_1
X_8437_ _3302_ _3322_ _3868_ _3331_ vssd1 vssd1 vccd1 vccd1 _3890_ sky130_fd_sc_hd__a31o_1
X_5649_ net61 _1526_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__xnor2_1
X_8368_ net81 _2240_ vssd1 vssd1 vccd1 vccd1 _3830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7319_ allocation.game.controller.init_module.delay_counter\[21\] _2967_ net123 vssd1
+ vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9356__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8299_ _3593_ _3751_ _3765_ net201 allocation.game.controller.drawBlock.y_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_5_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4526__X _0464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4951_ _0874_ _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__nand2_1
X_4882_ _0739_ _0762_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__nor2_2
X_7670_ _3213_ _3231_ vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__xor2_1
XANTENNA__4651__A_N allocation.game.controller.drawBlock.y_end\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6621_ allocation.game.cactusMove.count\[15\] allocation.game.cactusMove.count\[16\]
+ _2486_ allocation.game.cactusMove.count\[17\] vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__a31o_1
XANTENNA__9229__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9340_ clknet_leaf_3_clk allocation.game.collides net193 vssd1 vssd1 vccd1 vccd1
+ allocation.game.scoreCounter.col sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6552_ net468 _2441_ net90 vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6483_ allocation.game.scoreCounter.clock_div.counter\[4\] allocation.game.scoreCounter.clock_div.counter\[5\]
+ _2397_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__and3_1
X_5503_ _0795_ _0803_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__nor2_1
X_9271_ clknet_leaf_2_clk _0050_ net181 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9379__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8222_ _3033_ _3707_ _3708_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5434_ _1336_ _1358_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__xnor2_1
X_8153_ _0671_ _3639_ _3650_ allocation.game.controller.state\[7\] vssd1 vssd1 vccd1
+ vccd1 _3651_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7104_ _2809_ _2815_ _2816_ _2756_ vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_39_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5365_ _1283_ _1287_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5296_ _1161_ _1163_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__xnor2_1
X_8084_ net281 _3017_ _3467_ vssd1 vssd1 vccd1 vccd1 _3590_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_39_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7035_ _0417_ net4 vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_48_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8986_ _4432_ _4434_ _4430_ vssd1 vssd1 vccd1 vccd1 _4435_ sky130_fd_sc_hd__a21bo_1
X_7937_ allocation.game.controller.init_module.wr _3457_ _2926_ vssd1 vssd1 vccd1
+ vccd1 _0321_ sky130_fd_sc_hd__o21ba_1
XANTENNA__7657__X _3219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7868_ allocation.game.controller.drawBlock.state\[3\] net108 vssd1 vssd1 vccd1 vccd1
+ _3410_ sky130_fd_sc_hd__nor2_1
XANTENNA__7376__Y _3008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6819_ allocation.game.cactus2size.clock_div_inst0.counter\[0\] allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ allocation.game.cactus2size.clock_div_inst0.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2621_ sky130_fd_sc_hd__a21oi_1
X_7799_ _2861_ _3355_ vssd1 vssd1 vccd1 vccd1 _3361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9469_ clknet_leaf_8_clk _0376_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_end\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8648__B net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5353__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7727__B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5150_ _1071_ _1073_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__nor2_1
X_5081_ _0956_ _0961_ _1004_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6094__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8840_ net38 _4279_ _4289_ vssd1 vssd1 vccd1 vccd1 _4290_ sky130_fd_sc_hd__o21a_1
XANTENNA__9051__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5983_ _0778_ _0895_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__nor2_1
X_8771_ net40 _4220_ vssd1 vssd1 vccd1 vccd1 _4221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4934_ _0792_ _0817_ _0815_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__a21oi_1
X_7722_ net42 _3274_ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4865_ _0788_ _0789_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_9_clk_X clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7653_ allocation.game.lcdOutput.framebufferIndex\[9\] _3193_ _3204_ _3207_ _3203_
+ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__a41o_1
X_6604_ allocation.game.cactusMove.count\[10\] allocation.game.cactusMove.count\[11\]
+ _2477_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__and3_1
X_4796_ _0718_ _0719_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__nor2_1
X_7584_ net374 allocation.game.cactus2size.lfsr1\[1\] vssd1 vssd1 vccd1 vccd1 _3164_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9323_ clknet_leaf_6_clk _0106_ net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5760__A1 _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6535_ net475 _2430_ net90 vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7419__B1_N allocation.game.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9254_ clknet_leaf_0_clk _0075_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_8205_ _2377_ _3694_ _2379_ vssd1 vssd1 vccd1 vccd1 _3695_ sky130_fd_sc_hd__o21a_1
X_6466_ net234 net421 net232 vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6397_ allocation.game.scoreCounter.col _2315_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__or2_2
X_9185_ clknet_leaf_15_clk net328 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataShift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5417_ _1338_ _1340_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2_1
X_8136_ net239 _3634_ _3635_ _3631_ _3632_ vssd1 vssd1 vccd1 vccd1 _3636_ sky130_fd_sc_hd__a311o_1
X_5348_ _1217_ _1219_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_7_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8067_ net263 net136 _3479_ vssd1 vssd1 vccd1 vccd1 _3575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7018_ allocation.game.scoreCounter.bcd_tens\[5\] allocation.game.scoreCounter.bcd_tens\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__nor2_1
X_5279_ _1203_ _1202_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4804__X _0729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8969_ net129 _2253_ _2256_ net131 _4417_ vssd1 vssd1 vccd1 vccd1 _4418_ sky130_fd_sc_hd__o221a_1
XFILLER_0_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8394__A allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9074__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload7_A clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7738__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4650_ allocation.game.controller.drawBlock.y_start\[5\] allocation.game.controller.drawBlock.y_end\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4581_ _0498_ _0500_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__nand2_1
X_6320_ net259 _2240_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__nand2_1
X_6251_ allocation.game.controller.drawBlock.counter\[16\] _2175_ vssd1 vssd1 vccd1
+ vccd1 _2176_ sky130_fd_sc_hd__nor2_1
X_5202_ net73 _1070_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6182_ _2016_ _2106_ _2015_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9417__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5133_ _1011_ _1013_ _1056_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _0987_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__or2_1
X_8823_ net115 _3872_ net58 _3309_ vssd1 vssd1 vccd1 vccd1 _4273_ sky130_fd_sc_hd__or4b_1
XANTENNA__6758__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8754_ _4202_ _4204_ _4195_ vssd1 vssd1 vccd1 vccd1 _4205_ sky130_fd_sc_hd__a21o_1
X_5966_ _1886_ _1887_ _1889_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__nand3_1
X_4917_ _0797_ _0841_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__or2_2
XANTENNA__4784__A2 _0708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5897_ net103 net102 vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__nor2_1
XANTENNA__5981__A1 _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7705_ _3257_ _3265_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__nand2_1
X_8685_ _3208_ _3618_ _4129_ _4135_ vssd1 vssd1 vccd1 vccd1 _4136_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5718__D1 net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4848_ _0754_ _0772_ _0751_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__a21o_1
X_7636_ net125 allocation.game.lcdOutput.framebufferIndex\[11\] _3187_ _3195_ _3197_
+ vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_8_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4779_ _0582_ _0600_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__xnor2_2
X_7567_ allocation.game.lcdOutput.tft.spi.dataShift\[0\] allocation.game.lcdOutput.tft.spi.dataShift\[1\]
+ allocation.game.lcdOutput.tft.spi.dataShift\[2\] allocation.game.lcdOutput.tft.spi.dataShift\[3\]
+ allocation.game.lcdOutput.tft.spi.counter\[2\] allocation.game.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__mux4_1
X_9306_ clknet_leaf_21_clk _0079_ net189 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4800__A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7498_ net356 _0233_ _3109_ _3111_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__o22a_1
X_6518_ allocation.game.dinoJump.dinoDelay\[4\] _2419_ _2414_ vssd1 vssd1 vccd1 vccd1
+ _2422_ sky130_fd_sc_hd__o21ai_1
X_6449_ _2362_ _2367_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__nor2_1
X_9237_ clknet_leaf_22_clk _0021_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9168_ clknet_leaf_15_clk _0230_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9097__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8119_ _0616_ _3619_ vssd1 vssd1 vccd1 vccd1 _3620_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9059__RESET_B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9099_ clknet_leaf_14_clk _0195_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5631__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout47_X net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9195__D _0401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7740__B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9013__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6372__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5820_ _0896_ _1744_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_33_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5751_ _0819_ _1669_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5963__A1 _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4702_ net222 allocation.game.cactusMove.x_dist\[6\] vssd1 vssd1 vccd1 vccd1 _0629_
+ sky130_fd_sc_hd__nand2_1
X_8470_ _3922_ net34 _3359_ vssd1 vssd1 vccd1 vccd1 _3923_ sky130_fd_sc_hd__or3b_1
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5682_ _1576_ _1604_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__xnor2_1
X_7421_ _3023_ _3037_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4633_ allocation.game.controller.drawBlock.x_end\[0\] allocation.game.controller.drawBlock.x_start\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4564_ _0492_ _0501_ _0491_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__a21o_1
X_7352_ allocation.game.lcdOutput.tft.remainingDelayTicks\[14\] allocation.game.lcdOutput.tft.remainingDelayTicks\[13\]
+ _2991_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__or3_1
X_7283_ allocation.game.controller.init_module.delay_counter\[8\] _2942_ _2944_ vssd1
+ vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6303_ allocation.game.controller.drawBlock.counter\[19\] _2170_ _2227_ _2169_ vssd1
+ vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6234_ _1227_ _2131_ _1173_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__a21o_1
X_4495_ allocation.game.controller.drawBlock.counter\[20\] vssd1 vssd1 vccd1 vccd1
+ _0435_ sky130_fd_sc_hd__inv_2
X_9022_ net254 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8968__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6165_ net110 _0894_ _2081_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5451__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5116_ _1039_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__xnor2_1
X_6096_ _1987_ _1989_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__xnor2_1
X_5047_ _0931_ _0966_ _0967_ _0971_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6998_ allocation.game.bcd_ones\[0\] allocation.game.bcd_ones\[2\] vssd1 vssd1 vccd1
+ vccd1 _2735_ sky130_fd_sc_hd__xnor2_1
X_8806_ _3540_ _3760_ _4255_ vssd1 vssd1 vccd1 vccd1 _4256_ sky130_fd_sc_hd__a21bo_1
X_5949_ _1871_ _1872_ _1873_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__nand3_1
X_8737_ _4180_ _4187_ vssd1 vssd1 vccd1 vccd1 _4188_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8668_ _4096_ _4116_ _4117_ _4118_ vssd1 vssd1 vccd1 vccd1 _4119_ sky130_fd_sc_hd__or4b_1
XANTENNA__4801__Y _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7619_ allocation.game.lcdOutput.framebufferIndex\[16\] _2843_ _3180_ vssd1 vssd1
+ vccd1 vccd1 _3181_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8599_ net47 _4026_ vssd1 vssd1 vccd1 vccd1 _4050_ sky130_fd_sc_hd__nand2_1
XANTENNA__7841__A _3393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7092__C1 _0417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9112__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5945__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7934__A2 _3410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7735__B net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9262__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7970_ _3482_ vssd1 vssd1 vccd1 vccd1 _3483_ sky130_fd_sc_hd__inv_2
X_6921_ allocation.game.cactusDist.clock_div_inst0.counter\[7\] allocation.game.cactusDist.clock_div_inst0.counter\[8\]
+ _2685_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6852_ allocation.game.cactusDist.clock_div_inst1.counter\[1\] allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__or2_1
X_5803_ _1720_ _1727_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8522_ net58 _3337_ _3864_ _3872_ vssd1 vssd1 vccd1 vccd1 _3974_ sky130_fd_sc_hd__or4_1
X_6783_ _0448_ _2594_ _2597_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__a21oi_1
X_5734_ _1606_ _1607_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5665_ _1588_ _1589_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__nand2b_1
X_8453_ _3288_ _3869_ _3905_ _3344_ vssd1 vssd1 vccd1 vccd1 _3906_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout211_A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4616_ _0544_ _0545_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__nand2b_2
X_8384_ allocation.game.controller.v\[1\] allocation.game.controller.v\[0\] vssd1
+ vssd1 vccd1 vccd1 _3844_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7404_ _3001_ _3024_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__or2_1
X_7335_ _0436_ _2975_ _2980_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__o21ai_1
X_5596_ _1511_ _1513_ _1519_ _1520_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4547_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4478_ allocation.game.cactusMove.cactusMovement vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__inv_2
X_7266_ net420 _2931_ net122 vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__o21ai_1
X_7197_ allocation.game.dinoJump.count\[1\] allocation.game.dinoJump.count\[0\] allocation.game.dinoJump.count\[5\]
+ allocation.game.dinoJump.count\[4\] vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__and4_1
X_6217_ _1175_ _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__xnor2_1
X_9005_ _4450_ _4452_ _4453_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__and3_1
X_6148_ _0741_ _0895_ _2072_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__or3b_1
XANTENNA__9135__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6079_ _1965_ _2003_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9285__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8877__B1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7852__A1 allocation.game.controller.drawBlock.state\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5615__B1 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8801__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5091__A1 _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_14_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5450_ net61 _1373_ _1372_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5381_ net64 _1255_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7120_ _2828_ _2829_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7051_ allocation.game.controller.drawBlock.idx\[2\] allocation.game.controller.drawBlock.idx\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__nand2b_1
Xfanout219 net220 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
Xfanout208 net215 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
X_6002_ _1883_ _1925_ _1926_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__nand3_1
X_7953_ allocation.game.controller.state\[2\] allocation.game.controller.state\[7\]
+ _3466_ vssd1 vssd1 vccd1 vccd1 _3467_ sky130_fd_sc_hd__or3b_1
X_6904_ allocation.game.cactusDist.clock_div_inst0.counter\[1\] allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ allocation.game.cactusDist.clock_div_inst0.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2678_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout259_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7884_ _3420_ vssd1 vssd1 vccd1 vccd1 _3421_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout161_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6835_ allocation.game.cactus2size.clock_div_inst0.counter\[7\] _2629_ _2631_ vssd1
+ vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_18_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6766_ net334 _2583_ net154 vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5717_ _1639_ _1641_ _0911_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8505_ net132 net130 net126 vssd1 vssd1 vccd1 vccd1 _3957_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9485_ clknet_leaf_10_clk allocation.game.cactusMove.n_pixel\[5\] net202 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.pixel\[5\] sky130_fd_sc_hd__dfrtp_1
X_6697_ net158 _2539_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5648_ net61 _1571_ _1570_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__a21bo_1
X_8436_ _3888_ vssd1 vssd1 vccd1 vccd1 _3889_ sky130_fd_sc_hd__inv_2
X_8367_ _3479_ _3826_ _3828_ net242 vssd1 vssd1 vccd1 vccd1 _3829_ sky130_fd_sc_hd__o31a_1
XANTENNA__8487__A _3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5579_ _1502_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7318_ net123 _2966_ _2967_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__nor3_1
X_8298_ net281 _3752_ _3754_ _3764_ vssd1 vssd1 vccd1 vccd1 _3765_ sky130_fd_sc_hd__or4_1
XANTENNA__8087__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5904__A _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7249_ allocation.game.dinoJump.dinoMovement _0423_ _0529_ net278 _2919_ vssd1 vssd1
+ vccd1 vccd1 _2920_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout74_A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4807__X _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8653__C net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8397__A allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9300__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9005__B _4452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9021__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4950_ _0823_ _0873_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4881_ net71 _0802_ _0795_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__mux2_2
X_6620_ allocation.game.cactusMove.count\[17\] allocation.game.cactusMove.count\[16\]
+ _2487_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_41_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6551_ allocation.game.dinoJump.dinoDelay\[15\] allocation.game.dinoJump.dinoDelay\[16\]
+ _2439_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5502_ _0725_ _0820_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6482_ allocation.game.scoreCounter.clock_div.counter\[3\] _2396_ vssd1 vssd1 vccd1
+ vccd1 _2397_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9270_ clknet_leaf_2_clk _0049_ net177 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_8221_ _3019_ _3032_ _3001_ vssd1 vssd1 vccd1 vccd1 _3708_ sky130_fd_sc_hd__a21o_1
X_5433_ _1305_ _1357_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__nor2_1
XANTENNA__8069__B2 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8069__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8152_ net89 _3639_ vssd1 vssd1 vccd1 vccd1 _3650_ sky130_fd_sc_hd__nand2_1
X_5364_ _1235_ _1288_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7103_ allocation.game.controller.drawBlock.x_start\[7\] _2772_ _2777_ allocation.game.controller.drawBlock.x_end\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8083_ allocation.game.controller.drawBlock.y_start\[7\] net197 _3584_ _3589_ vssd1
+ vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_39_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5295_ _1217_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__nand2_1
X_7034_ _2755_ allocation.game.lcdOutput.tft.spi.tft_dc net4 vssd1 vssd1 vccd1 vccd1
+ net29 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8985_ _0657_ net52 _4431_ _4433_ vssd1 vssd1 vccd1 vccd1 _4434_ sky130_fd_sc_hd__o31a_1
X_7936_ allocation.game.controller.init_module.state\[0\] allocation.game.controller.init_module.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3457_ sky130_fd_sc_hd__and2b_1
X_7867_ allocation.game.controller.drawBlock.state\[2\] _3400_ _3402_ vssd1 vssd1
+ vccd1 vccd1 _3409_ sky130_fd_sc_hd__a21o_2
XFILLER_0_33_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6818_ net156 _2614_ _2620_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__and3_1
X_7798_ net35 _3359_ net39 vssd1 vssd1 vccd1 vccd1 _3360_ sky130_fd_sc_hd__o21ai_2
XANTENNA__7752__B1 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6749_ _2573_ _2574_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9323__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9468_ clknet_leaf_11_clk _0375_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_end\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8419_ net66 _3370_ vssd1 vssd1 vccd1 vccd1 _3872_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8010__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9399_ clknet_leaf_17_clk _0309_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8783__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8680__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7743__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8299__B2 allocation.game.controller.drawBlock.y_end\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9016__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5080_ _0956_ _0961_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5982_ net80 _1906_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6662__X _2516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8770_ net264 _4213_ vssd1 vssd1 vccd1 vccd1 _4220_ sky130_fd_sc_hd__xnor2_1
X_4933_ _0834_ _0841_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__nor2_1
X_7721_ _3282_ vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9106__RESET_B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4864_ _0786_ _0787_ _0773_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9346__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7652_ allocation.game.lcdOutput.framebufferIndex\[8\] _3204_ _3213_ vssd1 vssd1
+ vccd1 vccd1 _3214_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6603_ allocation.game.cactusMove.count\[10\] _2477_ _2479_ vssd1 vssd1 vccd1 vccd1
+ allocation.game.cactusMove.n_count\[10\] sky130_fd_sc_hd__o21a_1
X_4795_ _0718_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__and2_2
XFILLER_0_6_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7583_ net374 _2619_ _3014_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__mux2_1
X_9322_ clknet_leaf_6_clk _0129_ net173 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout124_A _0899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6534_ allocation.game.dinoJump.dinoDelay\[9\] allocation.game.dinoJump.dinoDelay\[10\]
+ _2428_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6465_ net237 net100 _2383_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9253_ clknet_leaf_1_clk _0074_ net169 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_8204_ _3692_ _3693_ vssd1 vssd1 vccd1 vccd1 _3694_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5454__A _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5416_ _1338_ _1340_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__or2_1
X_9184_ clknet_leaf_15_clk net347 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataShift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_6396_ _2316_ _2317_ allocation.game.scoreCounter.clock_div.slow_clk vssd1 vssd1
+ vccd1 vccd1 _2319_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_7_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8135_ net224 _0612_ net223 vssd1 vssd1 vccd1 vccd1 _3635_ sky130_fd_sc_hd__a21o_1
X_5347_ _1260_ _1263_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_7_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8765__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8066_ _3571_ _3572_ vssd1 vssd1 vccd1 vccd1 _3574_ sky130_fd_sc_hd__or2_1
X_5278_ _0834_ _1201_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__xnor2_1
X_7017_ _0450_ _0451_ allocation.game.bcd_ones\[2\] _2745_ _2747_ vssd1 vssd1 vccd1
+ vccd1 net18 sky130_fd_sc_hd__a311o_1
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8968_ net131 _2256_ _3312_ _4416_ vssd1 vssd1 vccd1 vccd1 _4417_ sky130_fd_sc_hd__a22o_1
X_7919_ net95 _3444_ _3445_ net109 allocation.game.controller.drawBlock.counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8899_ _4215_ _4348_ vssd1 vssd1 vccd1 vccd1 _4349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7844__A _2973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8675__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9219__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9369__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4580_ net235 _0515_ _0516_ net233 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoY\[5\]
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__5274__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6250_ _2114_ _2115_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__xnor2_1
XANTENNA__8692__A1 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5201_ _1124_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_36_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6181_ _2041_ _2105_ _2040_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5132_ _1011_ _1013_ _1056_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__o21a_1
Xclkbuf_1_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9514__299 vssd1 vssd1 vccd1 vccd1 _9514__299/HI net299 sky130_fd_sc_hd__conb_1
XFILLER_0_23_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5063_ _0986_ _0810_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__and2b_1
X_8822_ net258 _4245_ _4271_ vssd1 vssd1 vccd1 vccd1 _4272_ sky130_fd_sc_hd__a21o_1
X_8753_ _3219_ _4179_ _4197_ _4203_ _4191_ vssd1 vssd1 vccd1 vccd1 _4204_ sky130_fd_sc_hd__o311a_1
X_5965_ _1886_ _1887_ _1889_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__and3_1
X_4916_ _0728_ net79 vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__nor2_2
XANTENNA__5981__A2 _0729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7704_ _3257_ _3265_ vssd1 vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__and2_1
X_8684_ net76 _4123_ _4134_ vssd1 vssd1 vccd1 vccd1 _4135_ sky130_fd_sc_hd__o21ai_1
X_5896_ _1776_ _1818_ _1820_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__and3_1
X_4847_ _0766_ _0771_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__xnor2_4
XANTENNA__5718__C1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7635_ _3196_ net125 _3185_ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7566_ net353 allocation.game.lcdOutput.tft.spi.dataDc _2526_ vssd1 vssd1 vccd1 vccd1
+ _0253_ sky130_fd_sc_hd__mux2_1
X_4778_ _0585_ _0599_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__xnor2_4
X_9305_ clknet_leaf_22_clk _0078_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4800__B _0722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7497_ _3110_ net53 _3071_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__nand3b_1
X_6517_ allocation.game.dinoJump.dinoDelay\[3\] allocation.game.dinoJump.dinoDelay\[4\]
+ _2417_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__and3_1
X_6448_ net147 _2367_ _2369_ allocation.game.scoreCounter.bcd_tens\[5\] vssd1 vssd1
+ vccd1 vccd1 _0017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9236_ clknet_leaf_22_clk _0033_ net178 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6379_ net270 _2300_ _2302_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__o21ai_1
X_9167_ clknet_leaf_15_clk _0229_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8118_ net225 _0613_ vssd1 vssd1 vccd1 vccd1 _3619_ sky130_fd_sc_hd__and2_1
X_9098_ clknet_leaf_13_clk _0194_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_8049_ _3555_ _3557_ net135 vssd1 vssd1 vccd1 vccd1 _3558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4534__Y _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9041__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5750_ _1671_ _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__nand2_1
XANTENNA__5963__A2 _0729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4701_ net484 net238 _0609_ _0628_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a31o_1
X_5681_ _1599_ _1600_ _1602_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__o21ba_1
X_4632_ allocation.game.controller.drawBlock.x_start\[1\] allocation.game.controller.drawBlock.x_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__and2b_1
X_7420_ _3034_ _3038_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9472__Q allocation.game.controller.drawBlock.y_end\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4563_ _0498_ _0500_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__or2_1
X_7351_ allocation.game.lcdOutput.tft.remainingDelayTicks\[12\] _2990_ vssd1 vssd1
+ vccd1 vccd1 _2991_ sky130_fd_sc_hd__or2_1
X_7282_ allocation.game.controller.init_module.delay_counter\[8\] _2942_ _2927_ vssd1
+ vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6302_ allocation.game.controller.drawBlock.counter\[18\] _2172_ _2226_ _2171_ vssd1
+ vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__o211a_1
X_4494_ allocation.game.controller.drawBlock.counter\[19\] vssd1 vssd1 vccd1 vccd1
+ _0434_ sky130_fd_sc_hd__inv_2
X_6233_ _1119_ _2133_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_1_0__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7931__B _3409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9021_ net255 vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6164_ _0712_ _0894_ _2067_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__and3_1
X_5115_ _0841_ _0980_ _0983_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__or3_1
X_6095_ _1946_ _2019_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout191_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5046_ _0969_ _0970_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__and2b_1
XANTENNA__7378__B _3008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6997_ allocation.game.bcd_ones\[1\] allocation.game.bcd_ones\[3\] vssd1 vssd1 vccd1
+ vccd1 _2734_ sky130_fd_sc_hd__or2_1
X_8805_ net266 _4242_ vssd1 vssd1 vccd1 vccd1 _4255_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout244_X net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5948_ _1825_ _1870_ _1869_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__a21o_1
X_8736_ net121 _4179_ vssd1 vssd1 vccd1 vccd1 _4187_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8667_ net52 _3603_ vssd1 vssd1 vccd1 vccd1 _4118_ sky130_fd_sc_hd__xnor2_1
X_5879_ _0896_ _1695_ _1694_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__a21oi_1
X_7618_ allocation.game.lcdOutput.framebufferIndex\[16\] allocation.game.lcdOutput.framebufferIndex\[15\]
+ net125 allocation.game.lcdOutput.framebufferIndex\[13\] vssd1 vssd1 vccd1 vccd1
+ _3180_ sky130_fd_sc_hd__nand4_2
X_8598_ _4044_ _4048_ _4043_ vssd1 vssd1 vccd1 vccd1 _4049_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4530__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9064__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7549_ _3043_ _3149_ vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__nand2_1
XANTENNA__8656__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9219_ clknet_leaf_22_clk _0045_ net166 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7919__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9407__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5552__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5271__B _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6920_ allocation.game.cactusDist.clock_div_inst0.counter\[7\] _2685_ allocation.game.cactusDist.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9467__Q allocation.game.controller.drawBlock.y_end\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6851_ net358 _2639_ _2641_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__a21oi_1
X_5802_ _1720_ _1725_ _1726_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8521_ net114 _3972_ vssd1 vssd1 vccd1 vccd1 _3973_ sky130_fd_sc_hd__and2_1
X_6782_ net158 _2596_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__or2_1
XANTENNA__9087__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _1651_ _1655_ _1656_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__a21bo_1
X_5664_ _1121_ _1579_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__xor2_1
X_8452_ _3289_ _3321_ _3867_ _3904_ vssd1 vssd1 vccd1 vccd1 _3905_ sky130_fd_sc_hd__o31a_1
XFILLER_0_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8383_ allocation.game.controller.v\[1\] net84 vssd1 vssd1 vccd1 vccd1 _3843_ sky130_fd_sc_hd__and2b_1
X_4615_ allocation.game.controller.drawBlock.x_end\[7\] allocation.game.controller.drawBlock.x_start\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7403_ _3001_ _3024_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__nor2_1
X_5595_ _1466_ _1518_ _1517_ _1490_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_13_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4546_ allocation.game.controller.v\[5\] net265 vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7334_ _2977_ _2979_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4477_ net236 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7265_ allocation.game.controller.init_module.delay_counter\[2\] allocation.game.controller.init_module.delay_counter\[1\]
+ _2929_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__and3_1
XANTENNA__5462__A _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7196_ allocation.game.dinoJump.count\[3\] allocation.game.dinoJump.count\[2\] allocation.game.dinoJump.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__and3_1
X_6216_ _0793_ net71 _0802_ _0794_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9004_ _0462_ net216 _3272_ vssd1 vssd1 vccd1 vccd1 _4453_ sky130_fd_sc_hd__and3_1
X_6147_ _2070_ _2071_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__and2_1
XANTENNA__8810__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6078_ _1962_ _1964_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__or2_1
X_5029_ _0946_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_0_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8719_ net46 _4165_ _4169_ vssd1 vssd1 vccd1 vccd1 _4170_ sky130_fd_sc_hd__or3_1
XANTENNA__8877__A1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5457__A1_N _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5615__A1 _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7746__B net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9019__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8858__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5380_ net64 _1304_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_4
X_7050_ allocation.game.controller.drawBlock.idx\[4\] _2769_ vssd1 vssd1 vccd1 vccd1
+ _2770_ sky130_fd_sc_hd__or2_1
XANTENNA__7843__A2 _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6001_ _1879_ _1880_ _1882_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__a21o_1
X_7952_ net243 net239 _3465_ vssd1 vssd1 vccd1 vccd1 _3466_ sky130_fd_sc_hd__or3_1
X_6903_ allocation.game.cactusDist.clock_div_inst0.counter\[1\] allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ allocation.game.cactusDist.clock_div_inst0.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2677_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7883_ allocation.game.controller.drawBlock.counter\[4\] allocation.game.controller.drawBlock.counter\[5\]
+ _3415_ vssd1 vssd1 vccd1 vccd1 _3420_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_18_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout154_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6834_ allocation.game.cactus2size.clock_div_inst0.counter\[7\] _2629_ net160 vssd1
+ vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_18_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6765_ _2583_ _2584_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5716_ _0914_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__xnor2_1
X_9484_ clknet_leaf_10_clk allocation.game.cactusMove.n_pixel\[4\] net202 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.pixel\[4\] sky130_fd_sc_hd__dfrtp_1
X_8504_ _3947_ _3948_ _3955_ vssd1 vssd1 vccd1 vccd1 _3956_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8435_ _3331_ _3887_ vssd1 vssd1 vccd1 vccd1 _3888_ sky130_fd_sc_hd__nand2_1
X_6696_ _0447_ _2537_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5647_ _1570_ _1571_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8366_ net260 _3812_ _3827_ net140 vssd1 vssd1 vccd1 vccd1 _3828_ sky130_fd_sc_hd__o211a_1
X_5578_ _0773_ _1491_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__xor2_1
X_7317_ allocation.game.controller.init_module.delay_counter\[20\] allocation.game.controller.init_module.delay_counter\[19\]
+ _2963_ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__and3_1
X_8297_ net277 net163 _3556_ _3763_ vssd1 vssd1 vccd1 vccd1 _3764_ sky130_fd_sc_hd__a22o_1
XANTENNA__5904__B _0899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529_ net264 net261 vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__and2_2
X_7248_ _4458_ _0533_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__nor2_1
XANTENNA__9102__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7179_ net148 _2868_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9252__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8397__B allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6661__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4880_ _0800_ _0803_ _0795_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6550_ _2441_ _2442_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[15\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5501_ _1387_ _1425_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6481_ allocation.game.scoreCounter.clock_div.counter\[0\] allocation.game.scoreCounter.clock_div.counter\[2\]
+ allocation.game.scoreCounter.clock_div.counter\[1\] vssd1 vssd1 vccd1 vccd1 _2396_
+ sky130_fd_sc_hd__and3_1
XANTENNA__9125__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8220_ _2985_ _3706_ vssd1 vssd1 vccd1 vccd1 _3707_ sky130_fd_sc_hd__nand2_1
X_5432_ net64 _1304_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__nor2_1
X_8151_ _3637_ _3647_ vssd1 vssd1 vccd1 vccd1 _3649_ sky130_fd_sc_hd__nand2_1
X_5363_ _1234_ _1233_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7102_ allocation.game.controller.drawBlock.y_end\[7\] _2779_ _2787_ allocation.game.controller.drawBlock.y_start\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8082_ net259 net163 _3514_ _3588_ net281 vssd1 vssd1 vccd1 vccd1 _3589_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5294_ _1216_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__and2_1
XANTENNA__9275__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7033_ allocation.game.controller.init_module.wr allocation.game.controller.drawBlock.wr
+ net236 vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__mux2_1
XANTENNA__8844__A1_N net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8984_ _0652_ net57 vssd1 vssd1 vccd1 vccd1 _4433_ sky130_fd_sc_hd__nand2_1
X_7935_ _0435_ net109 _3455_ _3456_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__o31a_1
X_7866_ allocation.game.controller.drawBlock.idx\[4\] _3402_ vssd1 vssd1 vccd1 vccd1
+ _0299_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6817_ allocation.game.cactus2size.clock_div_inst0.counter\[0\] allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ _2619_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9536_ net317 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
X_7797_ _3311_ _3357_ vssd1 vssd1 vccd1 vccd1 _3359_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6748_ net450 _2571_ net153 vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6679_ _2526_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__inv_2
X_9467_ clknet_leaf_8_clk _0374_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_end\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9398_ clknet_leaf_17_clk _0308_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8418_ net66 net70 vssd1 vssd1 vccd1 vccd1 _3871_ sky130_fd_sc_hd__nor2_1
X_8349_ net263 _3795_ vssd1 vssd1 vccd1 vccd1 _3812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_13_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6491__B2 _0417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8768__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7991__A1 _3500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7743__A1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9148__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9405__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9298__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5809__A1 _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5981_ _0716_ _0729_ net83 vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__a21oi_1
X_4932_ _0842_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__and2_1
XANTENNA__6391__A _0462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7720_ net37 net35 vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__nor2_2
X_7651_ allocation.game.lcdOutput.framebufferIndex\[9\] net68 vssd1 vssd1 vccd1 vccd1
+ _3213_ sky130_fd_sc_hd__xnor2_2
X_6602_ allocation.game.cactusMove.count\[10\] _2477_ net145 vssd1 vssd1 vccd1 vccd1
+ _2479_ sky130_fd_sc_hd__a21oi_1
X_4863_ _0773_ _0786_ _0787_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__and3_1
X_4794_ _0561_ _0566_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__xnor2_1
X_7582_ net143 _3163_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9321_ clknet_leaf_6_clk _0128_ net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6533_ _2430_ _2431_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6464_ net237 _0626_ allocation.game.controller.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _2383_ sky130_fd_sc_hd__o21ai_1
X_9519__304 vssd1 vssd1 vccd1 vccd1 _9519__304/HI net304 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_31_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9252_ clknet_leaf_0_clk _0073_ net169 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8203_ net219 _2376_ vssd1 vssd1 vccd1 vccd1 _3693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5415_ _1293_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout117_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9183_ clknet_leaf_15_clk net341 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataShift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_6395_ allocation.game.scoreCounter.clock_div.slow_clk _2316_ vssd1 vssd1 vccd1 vccd1
+ _2318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8134_ _0612_ _2375_ vssd1 vssd1 vccd1 vccd1 _3634_ sky130_fd_sc_hd__nand2_1
X_5346_ _1267_ _1269_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_7_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8765__B net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8065_ _3571_ _3572_ vssd1 vssd1 vccd1 vccd1 _3573_ sky130_fd_sc_hd__nand2_1
X_5277_ _0797_ _1198_ _1200_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__a21o_1
X_7016_ _2740_ _2744_ _2747_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__or3_1
XFILLER_0_39_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8967_ allocation.game.cactusHeight2\[0\] allocation.game.cactusHeight2\[1\] _4415_
+ net133 vssd1 vssd1 vccd1 vccd1 _4416_ sky130_fd_sc_hd__a22o_1
XANTENNA__4814__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7918_ allocation.game.controller.drawBlock.counter\[15\] _3442_ vssd1 vssd1 vccd1
+ vccd1 _3445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8898_ _3811_ _4243_ _4345_ _3263_ _4216_ vssd1 vssd1 vccd1 vccd1 _4348_ sky130_fd_sc_hd__a221o_1
X_7849_ allocation.game.cactusHeight2\[5\] _2976_ _3394_ _3397_ vssd1 vssd1 vccd1
+ vccd1 _0292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9519_ net304 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XANTENNA__9440__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7844__B _3393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8021__A allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5200_ _1064_ _1122_ _1121_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_36_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6180_ _2102_ _2103_ _2048_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__a21o_1
X_5131_ _0798_ _1049_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5062_ _0810_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9313__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8821_ _4249_ _4267_ _4270_ _4263_ vssd1 vssd1 vccd1 vccd1 _4271_ sky130_fd_sc_hd__o22a_1
XANTENNA__7955__A1 allocation.game.collision.dinoY\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8752_ net69 _4188_ _4194_ vssd1 vssd1 vccd1 vccd1 _4203_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_17_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
X_7703_ allocation.game.lcdOutput.framebufferIndex\[4\] _3255_ vssd1 vssd1 vccd1 vccd1
+ _3265_ sky130_fd_sc_hd__or2_1
X_5964_ net110 net72 _1888_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__a21oi_1
X_4915_ _0837_ _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8683_ _4128_ _4131_ _4132_ _4133_ vssd1 vssd1 vccd1 vccd1 _4134_ sky130_fd_sc_hd__and4b_1
X_5895_ _1767_ _1773_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__xor2_2
XANTENNA__4921__X _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4846_ _0710_ _0770_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__nor2_4
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout234_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7634_ net125 _3180_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7565_ net398 _2527_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4777_ _0700_ _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__and2_2
X_9304_ clknet_leaf_22_clk _0077_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_6516_ _2419_ _2420_ net90 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7496_ allocation.game.lcdOutput.r_dino _3066_ _3068_ vssd1 vssd1 vccd1 vccd1 _3110_
+ sky130_fd_sc_hd__nor3_1
X_6447_ net147 _2360_ _2368_ _2369_ allocation.game.scoreCounter.bcd_tens\[6\] vssd1
+ vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9235_ clknet_leaf_22_clk _0032_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6378_ _2297_ _2298_ _2301_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__and3_1
X_9166_ clknet_leaf_15_clk _0228_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5329_ _1249_ _1251_ _1252_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__nand3_1
X_8117_ _3617_ vssd1 vssd1 vccd1 vccd1 _3618_ sky130_fd_sc_hd__inv_2
X_9097_ clknet_leaf_13_clk _0193_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_8048_ net265 _3542_ _3520_ vssd1 vssd1 vccd1 vccd1 _3557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9492__D _0392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9336__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9486__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9274__SET_B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4700_ net237 net113 vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _1576_ _1604_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4631_ _0559_ _0560_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__nand2b_1
X_4562_ net276 allocation.game.controller.v\[2\] vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__xnor2_2
X_7350_ allocation.game.lcdOutput.tft.remainingDelayTicks\[11\] allocation.game.lcdOutput.tft.remainingDelayTicks\[10\]
+ _2989_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7281_ _2942_ _2943_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6301_ allocation.game.controller.drawBlock.counter\[18\] _2172_ _2174_ _2225_ vssd1
+ vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__a211oi_1
X_4493_ allocation.game.controller.drawBlock.counter\[13\] vssd1 vssd1 vccd1 vccd1
+ _0433_ sky130_fd_sc_hd__inv_2
XANTENNA__8596__A _2516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_6_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
X_6232_ _1063_ _2134_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__xor2_1
X_9020_ net254 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6163_ _2085_ _2087_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__or2_1
X_5114_ _1037_ _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__nor2_1
X_6094_ net141 _0904_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__nor2_2
X_5045_ _0931_ _0968_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7640__A3 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8107__Y _3609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6996_ _0019_ _2733_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__nor2_1
X_8804_ net36 _4252_ vssd1 vssd1 vccd1 vccd1 _4254_ sky130_fd_sc_hd__nor2_1
X_5947_ _0770_ net124 vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__nor2_1
X_8735_ net120 _4183_ _4185_ net96 vssd1 vssd1 vccd1 vccd1 _4186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8666_ net59 _4098_ vssd1 vssd1 vccd1 vccd1 _4117_ sky130_fd_sc_hd__xnor2_1
XANTENNA__7675__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7617_ allocation.game.lcdOutput.framebufferIndex\[16\] allocation.game.lcdOutput.framebufferIndex\[15\]
+ net125 _0440_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__a31o_1
X_5878_ _1764_ _1802_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__and2b_1
X_4829_ _0751_ _0753_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8597_ net58 _3609_ _4045_ _4046_ _4047_ vssd1 vssd1 vccd1 vccd1 _4048_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4914__A1 _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7548_ _3040_ _3149_ net249 vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8656__A2 _3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7479_ _0430_ net250 vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__nand2_1
XANTENNA__9359__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9218_ clknet_leaf_0_clk _0044_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout97_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9149_ clknet_leaf_9_clk _0213_ net196 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.x_dist\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__8408__A2 _3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5890__A2 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7092__B2 allocation.game.controller.drawBlock.y_end\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6754__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7919__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1 allocation.game.sync0 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6850_ net358 _2639_ net156 vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4654__A_N allocation.game.controller.drawBlock.y_end\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5801_ _1674_ _1719_ net80 vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6781_ _0448_ _2594_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5732_ _1655_ _1656_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__xnor2_1
X_8520_ _3369_ _3892_ _3371_ vssd1 vssd1 vccd1 vccd1 _3972_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5663_ _1586_ _1587_ _1581_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__a21oi_1
X_8451_ _3322_ _3868_ _3290_ vssd1 vssd1 vccd1 vccd1 _3904_ sky130_fd_sc_hd__a21o_1
X_8382_ allocation.game.controller.v\[0\] _3842_ _3837_ vssd1 vssd1 vccd1 vccd1 _0381_
+ sky130_fd_sc_hd__o21ai_1
X_4614_ allocation.game.controller.drawBlock.x_start\[7\] allocation.game.controller.drawBlock.x_end\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5594_ _1490_ _1517_ _1518_ _1466_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7402_ allocation.game.lcdOutput.tft.state\[2\] net256 _3023_ allocation.game.lcdOutput.tft.spi.idle
+ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__or4b_2
X_4545_ net265 allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__and2b_1
X_7333_ _2973_ _2978_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7264_ _2931_ _2932_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__nor2_1
X_4476_ allocation.game.controller.drawBlock.x_end\[8\] vssd1 vssd1 vccd1 vccd1 _0416_
+ sky130_fd_sc_hd__inv_2
X_9003_ net35 _3274_ _4451_ net39 vssd1 vssd1 vccd1 vccd1 _4452_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7195_ net84 _2877_ _2879_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__and3_1
X_6215_ _1026_ _1032_ _1030_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6146_ _2019_ _2067_ _2069_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6077_ _1999_ _2001_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__nand2_1
X_5028_ _0871_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4806__B net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6979_ allocation.game.scoreCounter.clock_div.counter\[17\] _2721_ allocation.game.scoreCounter.clock_div.counter\[18\]
+ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__a21o_1
XANTENNA__9031__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8326__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4822__A _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8718_ _4095_ _4168_ vssd1 vssd1 vccd1 vccd1 _4169_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_7_clk_X clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8649_ net121 _4097_ vssd1 vssd1 vccd1 vccd1 _4100_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7837__A0 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5615__A2 _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7867__X _3409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5828__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5282__B _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6000_ _1863_ _1922_ _1923_ _1924_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__nor4_2
XANTENNA__7056__A1 allocation.game.controller.drawBlock.x_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9478__Q allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7951_ net242 allocation.game.controller.state\[0\] _2413_ vssd1 vssd1 vccd1 vccd1
+ _3465_ sky130_fd_sc_hd__or3_1
XANTENNA__9054__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7882_ net94 _3418_ _3419_ net108 allocation.game.controller.drawBlock.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__a32o_1
X_6902_ net155 _2673_ _2675_ _2676_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6833_ _2629_ _2630_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout147_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6764_ net466 _2582_ net154 vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5715_ net102 _0909_ _0910_ _0800_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__a211o_1
X_9483_ clknet_leaf_11_clk allocation.game.cactusMove.n_pixel\[3\] net202 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.pixel\[3\] sky130_fd_sc_hd__dfstp_1
X_6695_ net153 _2534_ _2537_ _2538_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__and4_1
X_8503_ _3883_ _3949_ _3951_ _3953_ _3954_ vssd1 vssd1 vccd1 vccd1 _3955_ sky130_fd_sc_hd__o32a_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5646_ _1521_ _1569_ _1568_ _1564_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__o211ai_1
X_8434_ _3200_ net68 _3297_ vssd1 vssd1 vccd1 vccd1 _3887_ sky130_fd_sc_hd__or3_1
X_8365_ net260 _3812_ vssd1 vssd1 vccd1 vccd1 _3827_ sky130_fd_sc_hd__nand2_1
X_5577_ _0831_ _1493_ _1501_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__a21bo_1
X_7316_ allocation.game.controller.init_module.delay_counter\[19\] _2963_ allocation.game.controller.init_module.delay_counter\[20\]
+ vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__a21oi_1
X_8296_ net134 _3757_ _3758_ _3762_ vssd1 vssd1 vccd1 vccd1 _3763_ sky130_fd_sc_hd__a31o_1
X_4528_ net275 _4458_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__and2_1
X_7247_ net275 allocation.game.dinoJump.next_dinoY\[2\] vssd1 vssd1 vccd1 vccd1 _2918_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7178_ allocation.game.dinoJump.count\[1\] allocation.game.dinoJump.count\[0\] allocation.game.dinoJump.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__and3_1
XANTENNA__5920__B _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4817__A _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6129_ _0715_ _0904_ _0908_ net141 vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_5_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9077__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5500_ _0731_ _1386_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__or2_1
X_6480_ allocation.game.scoreCounter.clock_div.counter\[19\] _2387_ _2394_ allocation.game.scoreCounter.clock_div.counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__o211a_1
XANTENNA__8710__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8710__B2 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5524__A1 _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5431_ net64 _1355_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__nand2_1
X_8150_ _3637_ _3647_ vssd1 vssd1 vccd1 vccd1 _3648_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5362_ _1284_ _1286_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7101_ _2809_ _2813_ _2814_ _2760_ vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__o31a_1
X_8081_ net259 net140 _3586_ _3587_ vssd1 vssd1 vccd1 vccd1 _3588_ sky130_fd_sc_hd__o22a_1
X_7032_ allocation.game.lcdOutput.tft.tft_reset net4 vssd1 vssd1 vccd1 vccd1 net30
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_39_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5293_ _1193_ _1213_ _1215_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8983_ _4149_ _4171_ _4431_ vssd1 vssd1 vccd1 vccd1 _4432_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout264_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7934_ allocation.game.controller.drawBlock.counter\[19\] _3410_ _3452_ allocation.game.controller.drawBlock.counter\[20\]
+ vssd1 vssd1 vccd1 vccd1 _3456_ sky130_fd_sc_hd__a31o_1
X_7865_ allocation.game.controller.drawBlock.idx\[3\] _3407_ _3408_ _3403_ vssd1 vssd1
+ vccd1 vccd1 _0298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7667__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5468__A _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8544__A4 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6816_ _2616_ _2617_ _2618_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__nor3_1
X_7796_ net42 _3356_ vssd1 vssd1 vccd1 vccd1 _3358_ sky130_fd_sc_hd__nand2_1
X_9535_ net316 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6747_ allocation.game.cactus1size.clock_div_inst0.counter\[5\] allocation.game.cactus1size.clock_div_inst0.counter\[6\]
+ _2569_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6678_ net422 _0431_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__nor2_4
XFILLER_0_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9466_ clknet_leaf_11_clk _0373_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_end\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5629_ _0728_ _0770_ _1066_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__o21ai_2
X_9397_ clknet_leaf_17_clk _0307_ net215 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_8417_ _3324_ _3868_ vssd1 vssd1 vccd1 vccd1 _3870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8348_ net266 net262 vssd1 vssd1 vccd1 vccd1 _3811_ sky130_fd_sc_hd__nor2_1
X_8279_ net137 _3472_ vssd1 vssd1 vccd1 vccd1 _3747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4834__X _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6762__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8940__B2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7593__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5980_ _1902_ _1903_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__xnor2_1
X_4931_ _0797_ _0834_ _0804_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__o21a_1
XANTENNA__6391__B _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5993__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4862_ _0780_ _0785_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__or2_1
X_7650_ _3193_ _3211_ vssd1 vssd1 vccd1 vccd1 _3212_ sky130_fd_sc_hd__xor2_1
X_6601_ _2477_ _2478_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9320_ clknet_leaf_6_clk _0127_ net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4793_ _0711_ _0563_ _0565_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__mux2_2
X_7581_ allocation.game.cactus1size.lfsr2\[1\] allocation.game.cactus1size.lfsr2\[0\]
+ allocation.game.cactus1size.clock_div_inst1.clk1 vssd1 vssd1 vccd1 vccd1 _3163_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8599__A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6532_ allocation.game.dinoJump.dinoDelay\[9\] _2428_ _2415_ vssd1 vssd1 vccd1 vccd1
+ _2431_ sky130_fd_sc_hd__o21ai_1
X_6463_ net239 _2380_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9242__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9251_ clknet_leaf_1_clk _0072_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_8202_ net222 allocation.game.cactusMove.pixel\[7\] _2311_ vssd1 vssd1 vccd1 vccd1
+ _3692_ sky130_fd_sc_hd__and3_1
X_9182_ clknet_leaf_15_clk net336 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataShift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_5414_ _1031_ _1292_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8133_ _3632_ vssd1 vssd1 vccd1 vccd1 _3633_ sky130_fd_sc_hd__inv_2
X_6394_ allocation.game.game.score\[3\] allocation.game.game.score\[2\] allocation.game.game.score\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__nor3_1
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5345_ _1246_ _1266_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_7_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8998__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8064_ _3531_ _3534_ _3543_ _3544_ vssd1 vssd1 vccd1 vccd1 _3572_ sky130_fd_sc_hd__a31o_1
X_5276_ _1197_ _1199_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__xnor2_4
XANTENNA__9392__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7015_ _0451_ _2737_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8966_ _0401_ allocation.game.cactusHeight2\[0\] allocation.game.cactusHeight2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _4415_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4814__B net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7917_ allocation.game.controller.drawBlock.counter\[15\] _3442_ vssd1 vssd1 vccd1
+ vccd1 _3444_ sky130_fd_sc_hd__or2_1
X_8897_ _4344_ _4346_ _4257_ _4343_ vssd1 vssd1 vccd1 vccd1 _4347_ sky130_fd_sc_hd__a211oi_1
X_7848_ net462 _2975_ _3396_ _3398_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__o211a_1
X_7779_ _3253_ net42 vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9518_ net303 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XANTENNA__8047__A_N net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9449_ clknet_leaf_18_clk _0356_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout82_X net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7588__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9115__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Left_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8913__A1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9265__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5130_ net62 _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5061_ _0809_ _0819_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__xor2_1
X_8820_ _4254_ _4269_ _4253_ vssd1 vssd1 vccd1 vccd1 _4270_ sky130_fd_sc_hd__o21ba_1
XANTENNA__7955__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8751_ _3228_ _4196_ _4198_ _4201_ vssd1 vssd1 vccd1 vccd1 _4202_ sky130_fd_sc_hd__a211o_1
X_5963_ _0722_ _0729_ net72 vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4914_ _0710_ _0799_ _0838_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__o21bai_1
XANTENNA__4634__B allocation.game.controller.drawBlock.x_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_7702_ _3239_ _3262_ vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5894_ _1772_ _1812_ _1817_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__nand3_1
X_8682_ _4125_ _4130_ net98 vssd1 vssd1 vccd1 vccd1 _4133_ sky130_fd_sc_hd__o21ai_1
X_4845_ _0758_ _0767_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_34_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7633_ _3187_ _3192_ vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4776_ _0596_ _0598_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__xnor2_4
X_7564_ _2527_ _3154_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__nor2_1
XANTENNA__5746__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9303_ clknet_leaf_22_clk _0089_ net180 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6515_ allocation.game.dinoJump.dinoDelay\[3\] _2417_ vssd1 vssd1 vccd1 vccd1 _2420_
+ sky130_fd_sc_hd__or2_1
X_7495_ net246 _3105_ _3108_ vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__o21ba_1
X_6446_ net234 _4455_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__nor2_2
XANTENNA__6143__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9234_ clknet_leaf_22_clk _0031_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6377_ net266 _2295_ _2300_ net271 vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__a22oi_1
X_9165_ clknet_leaf_16_clk _0227_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9096_ clknet_leaf_13_clk _0192_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_8116_ _0689_ _3616_ vssd1 vssd1 vccd1 vccd1 _3617_ sky130_fd_sc_hd__or2_2
X_5328_ _1249_ _1251_ _1252_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__a21o_1
X_8047_ net107 net241 vssd1 vssd1 vccd1 vccd1 _3556_ sky130_fd_sc_hd__and2b_1
X_5259_ _0842_ _1139_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_43_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7201__A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8949_ net75 _4395_ _4397_ vssd1 vssd1 vccd1 vccd1 _4398_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9288__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload5_A clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4630_ allocation.game.controller.drawBlock.x_end\[2\] allocation.game.controller.drawBlock.x_start\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__nand2b_1
XANTENNA__4470__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4561_ allocation.game.controller.v\[2\] net276 vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6300_ allocation.game.controller.drawBlock.counter\[17\] _2173_ _2176_ _2224_ vssd1
+ vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__a211o_1
X_7280_ net483 _2941_ net122 vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4492_ allocation.game.controller.drawBlock.counter\[11\] vssd1 vssd1 vccd1 vccd1
+ _0432_ sky130_fd_sc_hd__inv_2
X_6231_ _2135_ _2155_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6162_ _2076_ _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__or2_1
X_5113_ _1015_ _1036_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6093_ _0761_ _0894_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__nand2_1
X_5044_ _0924_ _0928_ _0926_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__o21a_1
XANTENNA__9430__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8803_ net38 _4250_ _4252_ net36 vssd1 vssd1 vccd1 vccd1 _4253_ sky130_fd_sc_hd__a22o_1
X_6995_ allocation.game.scoreCounter.clock_div.counter\[23\] _2730_ net386 vssd1 vssd1
+ vccd1 vccd1 _2733_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5946_ _1825_ _1869_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__nand3_1
X_8734_ net104 _4181_ vssd1 vssd1 vccd1 vccd1 _4185_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5877_ _1765_ _1801_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__and2b_1
X_8665_ _4097_ _4099_ _4115_ vssd1 vssd1 vccd1 vccd1 _4116_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4828_ _0746_ _0750_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__and2b_1
X_7616_ net125 allocation.game.lcdOutput.framebufferIndex\[11\] vssd1 vssd1 vccd1
+ vccd1 _3178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8596_ _2516_ net52 _4012_ vssd1 vssd1 vccd1 vccd1 _4047_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4759_ _0654_ _0685_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__nand2_1
X_7547_ net251 _3055_ _3039_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__mux2_1
X_7478_ _3048_ _3051_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__nand2_1
X_6429_ _2351_ _0421_ _2320_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__mux2_1
X_9217_ clknet_leaf_0_clk _0043_ net169 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4678__A1 _0417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9148_ clknet_leaf_10_clk _0212_ net196 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.x_dist\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_9079_ clknet_leaf_14_clk _0175_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9504__289 vssd1 vssd1 vccd1 vccd1 _9504__289/HI net289 sky130_fd_sc_hd__conb_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9303__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2 allocation.game.dinoJump.button vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5800_ _1723_ _1724_ _1722_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6780_ _2592_ _2594_ _2595_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5731_ _1578_ _1603_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5662_ _0784_ _1580_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__xnor2_1
X_8450_ _3877_ _3886_ _3902_ _3861_ vssd1 vssd1 vccd1 vccd1 _3903_ sky130_fd_sc_hd__a31o_1
X_8381_ _3840_ _3841_ vssd1 vssd1 vccd1 vccd1 _3842_ sky130_fd_sc_hd__nand2_2
X_4613_ allocation.game.controller.drawBlock.x_start\[8\] _0416_ vssd1 vssd1 vccd1
+ vccd1 _0543_ sky130_fd_sc_hd__nor2_1
X_5593_ _1439_ _1464_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__or2_1
X_7401_ _3021_ _3022_ allocation.game.lcdOutput.tft.state\[0\] _3018_ vssd1 vssd1
+ vccd1 vccd1 _3023_ sky130_fd_sc_hd__o211a_1
X_4544_ _4459_ _0481_ net235 vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__o21a_1
X_7332_ allocation.game.cactus1size.lfsr1\[0\] allocation.game.cactus1size.lfsr2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__xor2_2
X_7263_ net469 _2929_ net122 vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4475_ net219 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__inv_2
X_6214_ _1039_ _1040_ _1037_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__a21o_1
X_9002_ net131 _3312_ net45 net129 vssd1 vssd1 vccd1 vccd1 _4451_ sky130_fd_sc_hd__a211o_1
X_7194_ _2875_ _2878_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6145_ _2019_ _2067_ _2069_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__nand3_1
X_6076_ _1859_ _2000_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__nor2_1
X_5027_ _0950_ _0951_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__and2_1
XANTENNA__6282__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6978_ net390 _2721_ _2722_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_24_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8717_ _4141_ _4167_ vssd1 vssd1 vccd1 vccd1 _4168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5929_ _1849_ _1850_ _1853_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9326__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8648_ net121 net69 vssd1 vssd1 vccd1 vccd1 _4099_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8579_ _4025_ _4029_ _3996_ vssd1 vssd1 vccd1 vccd1 _4030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5934__A _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9476__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6328__A1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7950_ net243 net239 net281 vssd1 vssd1 vccd1 vccd1 _3464_ sky130_fd_sc_hd__or3_1
X_7881_ allocation.game.controller.drawBlock.counter\[4\] _3415_ vssd1 vssd1 vccd1
+ vccd1 _3419_ sky130_fd_sc_hd__or2_1
X_6901_ allocation.game.cactusDist.clock_div_inst0.counter\[1\] allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__nand2_1
XANTENNA__4771__A_N allocation.game.controller.drawBlock.y_start\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6832_ net482 _2627_ net156 vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9349__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6763_ allocation.game.cactus1size.clock_div_inst0.counter\[12\] _2582_ vssd1 vssd1
+ vccd1 vccd1 _2583_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9482_ clknet_leaf_11_clk allocation.game.cactusMove.n_pixel\[2\] net202 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.pixel\[2\] sky130_fd_sc_hd__dfrtp_1
X_5714_ _1635_ _1636_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__a21oi_1
X_6694_ allocation.game.cactus1size.clock_div_inst1.counter\[1\] allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ allocation.game.cactus1size.clock_div_inst1.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2538_ sky130_fd_sc_hd__a21o_1
X_8502_ _3327_ _3864_ net70 net117 vssd1 vssd1 vccd1 vccd1 _3954_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5645_ _1564_ _1568_ _1569_ _1521_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__a211o_1
X_8433_ _3277_ _3879_ _3885_ _3878_ vssd1 vssd1 vccd1 vccd1 _3886_ sky130_fd_sc_hd__or4b_1
XFILLER_0_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8364_ net136 _3824_ _3825_ vssd1 vssd1 vccd1 vccd1 _3826_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5576_ _1500_ _1499_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__nand2b_1
X_7315_ allocation.game.controller.init_module.delay_counter\[19\] _2963_ _2965_ vssd1
+ vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__o21a_1
X_8295_ _3759_ _3761_ net134 vssd1 vssd1 vccd1 vccd1 _3762_ sky130_fd_sc_hd__a21oi_1
X_4527_ _0461_ _0464_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7246_ net264 allocation.game.dinoJump.next_dinoY\[5\] vssd1 vssd1 vccd1 vccd1 _2917_
+ sky130_fd_sc_hd__or2_1
X_7177_ allocation.game.dinoJump.count\[1\] allocation.game.dinoJump.count\[0\] net148
+ allocation.game.dinoJump.count\[2\] vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6128_ _2043_ _2045_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_5_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _1970_ _1971_ _1967_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_29_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5430_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__and2_1
XANTENNA__5524__A2 _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5361_ _1283_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__nor2_1
X_8080_ _3569_ _3574_ _3585_ net136 vssd1 vssd1 vccd1 vccd1 _3587_ sky130_fd_sc_hd__a31o_1
X_7100_ allocation.game.controller.drawBlock.x_start\[6\] _2772_ _2777_ allocation.game.controller.drawBlock.x_end\[6\]
+ _2812_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__a221o_1
X_5292_ _1208_ _1211_ _1209_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8474__A1 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7031_ allocation.game.scoreCounter.bcd_tens\[6\] allocation.game.scoreCounter.bcd_tens\[3\]
+ _2752_ _0445_ _0446_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__o311a_1
XANTENNA__4918__A _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_X clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8982_ _0652_ _3219_ vssd1 vssd1 vccd1 vccd1 _4431_ sky130_fd_sc_hd__nor2_1
X_7933_ allocation.game.controller.drawBlock.counter\[19\] _3452_ _3454_ _3455_ vssd1
+ vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__o22a_1
X_7864_ _2762_ _2774_ _3400_ vssd1 vssd1 vccd1 vccd1 _3408_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7795_ net132 _3355_ vssd1 vssd1 vccd1 vccd1 _3357_ sky130_fd_sc_hd__or2_1
X_6815_ allocation.game.cactus2size.clock_div_inst0.counter\[11\] allocation.game.cactus2size.clock_div_inst0.counter\[10\]
+ allocation.game.cactus2size.clock_div_inst0.counter\[13\] allocation.game.cactus2size.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9534_ net315 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
X_6746_ _2571_ _2572_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6677_ net218 _2525_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_pixel\[8\]
+ sky130_fd_sc_hd__xnor2_1
X_9465_ clknet_leaf_1_clk _0372_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4667__A_N allocation.game.controller.drawBlock.y_end\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9396_ clknet_leaf_17_clk _0306_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_8416_ _3297_ _3866_ vssd1 vssd1 vccd1 vccd1 _3869_ sky130_fd_sc_hd__nor2_1
X_5628_ net65 _1508_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__xor2_1
X_8347_ net263 _3795_ vssd1 vssd1 vccd1 vccd1 _3810_ sky130_fd_sc_hd__and2_1
X_5559_ _0732_ _1483_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8278_ net279 _3483_ net136 vssd1 vssd1 vccd1 vccd1 _3746_ sky130_fd_sc_hd__mux2_1
X_7229_ allocation.game.dinoJump.count\[15\] allocation.game.dinoJump.count\[16\]
+ _2900_ allocation.game.dinoJump.count\[17\] vssd1 vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout72_A _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8768__A2 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5659__A _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8035__A allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9044__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6429__S _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9194__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _0834_ _0842_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__or2_1
X_4861_ _0780_ _0785_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__nand2_1
X_6600_ allocation.game.cactusMove.count\[9\] _2475_ net149 vssd1 vssd1 vccd1 vccd1
+ _2478_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7580_ _3161_ _3162_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__nor2_1
X_4792_ net83 _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6531_ allocation.game.dinoJump.dinoDelay\[9\] _2428_ vssd1 vssd1 vccd1 vccd1 _2430_
+ sky130_fd_sc_hd__and2_1
X_6462_ _2380_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8695__A1 net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9250_ clknet_leaf_1_clk _0071_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_8201_ _0692_ _3690_ net77 vssd1 vssd1 vccd1 vccd1 _3691_ sky130_fd_sc_hd__a21oi_1
X_9181_ clknet_leaf_15_clk net344 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataShift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6393_ allocation.game.game.score\[6\] allocation.game.game.score\[5\] vssd1 vssd1
+ vccd1 vccd1 _2316_ sky130_fd_sc_hd__nand2_2
XFILLER_0_3_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5413_ _0992_ _1337_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__or2_1
X_8132_ allocation.game.controller.state\[0\] net282 vssd1 vssd1 vccd1 vccd1 _3632_
+ sky130_fd_sc_hd__or2_1
X_5344_ _1213_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7950__C net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8063_ _3569_ _3570_ vssd1 vssd1 vccd1 vccd1 _3571_ sky130_fd_sc_hd__nand2_1
X_5275_ _1197_ _1199_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__and2b_1
XANTENNA__8998__A2 _3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7014_ allocation.game.bcd_ones\[0\] _2737_ _2746_ vssd1 vssd1 vccd1 vccd1 net16
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8965_ _4401_ _4404_ _4408_ _4413_ vssd1 vssd1 vccd1 vccd1 _4414_ sky130_fd_sc_hd__a31oi_1
X_7916_ _3442_ _3443_ allocation.game.controller.drawBlock.counter\[14\] net109 vssd1
+ vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a2bb2o_1
X_8896_ net35 _4345_ vssd1 vssd1 vccd1 vccd1 _4346_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout162_X net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7847_ allocation.game.cactusHeight2\[3\] _2976_ _3395_ _3397_ vssd1 vssd1 vccd1
+ vccd1 _0290_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ _3330_ _3339_ _3316_ vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9517_ net302 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XANTENNA__9067__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6729_ _2558_ _2560_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9448_ clknet_leaf_18_clk _0355_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9379_ clknet_leaf_10_clk _0289_ net196 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4829__Y _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8972__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4468__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5060_ _0983_ _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__or2_1
X_8750_ _3228_ _4196_ _4199_ _4200_ vssd1 vssd1 vccd1 vccd1 _4201_ sky130_fd_sc_hd__o22a_1
X_5962_ _1840_ _1885_ _1884_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__a21o_1
X_4913_ net88 _0764_ _0765_ _0771_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__a22o_2
X_7701_ _3239_ _3262_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__xor2_2
X_9525__310 vssd1 vssd1 vccd1 vccd1 _9525__310/HI net310 sky130_fd_sc_hd__conb_1
X_5893_ _1772_ _1812_ _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__and3_1
X_8681_ net120 _4127_ vssd1 vssd1 vccd1 vccd1 _4132_ sky130_fd_sc_hd__nand2_1
XANTENNA__8403__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4844_ _0758_ _0767_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__xor2_4
XFILLER_0_34_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7632_ allocation.game.lcdOutput.framebufferIndex\[10\] _3187_ _3193_ vssd1 vssd1
+ vccd1 vccd1 _3194_ sky130_fd_sc_hd__nand3_1
XANTENNA__4650__B allocation.game.controller.drawBlock.y_end\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4775_ _0594_ _0698_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__and3_4
X_7563_ allocation.game.lcdOutput.tft.spi.counter\[2\] _2526_ net415 vssd1 vssd1 vccd1
+ vccd1 _3154_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5746__B _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9302_ clknet_leaf_22_clk _0088_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6514_ allocation.game.dinoJump.dinoDelay\[3\] _2417_ vssd1 vssd1 vccd1 vccd1 _2419_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7494_ net246 _3106_ _3107_ _3020_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__a31o_1
X_9233_ clknet_leaf_22_clk _0030_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6445_ _2361_ _2367_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6376_ _2291_ _2299_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__or2_1
X_9164_ clknet_leaf_16_clk _0226_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_9095_ clknet_leaf_14_clk _0191_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8115_ _0688_ net121 vssd1 vssd1 vccd1 vccd1 _3616_ sky130_fd_sc_hd__and2b_1
X_5327_ _1202_ _1203_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__xor2_1
X_9532__314 vssd1 vssd1 vccd1 vccd1 _9532__314/HI net314 sky130_fd_sc_hd__conb_1
X_8046_ _0486_ _3554_ vssd1 vssd1 vccd1 vccd1 _3555_ sky130_fd_sc_hd__xnor2_1
X_5258_ _1027_ _1182_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__nor2_1
X_5189_ net62 _1113_ _1111_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8948_ net97 _3694_ vssd1 vssd1 vccd1 vccd1 _4397_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8356__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8879_ net266 _4308_ _4328_ vssd1 vssd1 vccd1 vccd1 _4329_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout35_A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6842__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
Xfanout180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
XANTENNA__9232__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9382__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4908__A0 _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4560_ net278 allocation.game.controller.v\[1\] _0497_ vssd1 vssd1 vccd1 vccd1 _0498_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4491_ net447 vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6230_ _2136_ _2154_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__xnor2_1
X_6161_ _2070_ _2073_ _2075_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__and3_1
X_5112_ _1015_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__and2_1
X_6092_ _2015_ _2016_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__and2b_1
XANTENNA__8822__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5043_ _0966_ _0967_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__nand2_1
XANTENNA__8050__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8802_ _4245_ _4251_ vssd1 vssd1 vccd1 vccd1 _4252_ sky130_fd_sc_hd__or2_1
X_6994_ net378 _2730_ _2732_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5945_ net87 _0903_ _1823_ _1824_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__a22o_1
X_8733_ net120 _4183_ vssd1 vssd1 vccd1 vccd1 _4184_ sky130_fd_sc_hd__nor2_1
X_5876_ _1796_ _1797_ _1800_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__a21o_1
X_8664_ _4097_ _4099_ _4100_ _4109_ _4114_ vssd1 vssd1 vccd1 vccd1 _4115_ sky130_fd_sc_hd__o221a_1
XANTENNA__8889__B2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8889__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4827_ _0751_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__inv_2
X_7615_ net232 allocation.game.game.score\[6\] net146 _2341_ vssd1 vssd1 vccd1 vccd1
+ _0279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8595_ net229 _3292_ _3863_ vssd1 vssd1 vccd1 vccd1 _4046_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7546_ _3039_ _3077_ _3150_ net252 vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4758_ net257 net164 vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4689_ allocation.game.cactusMove.pixel\[5\] _0613_ vssd1 vssd1 vccd1 vccd1 _0617_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_31_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7477_ net248 _3050_ _3083_ _3057_ _3051_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__a32o_1
XANTENNA__9105__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6428_ _2321_ _2350_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9216_ clknet_leaf_0_clk _0042_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_9147_ clknet_leaf_10_clk _0211_ net196 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.x_dist\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ net277 _2282_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9078_ clknet_leaf_14_clk _0174_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5627__A1 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8029_ allocation.game.controller.drawBlock.y_start\[4\] net197 _3537_ _3538_ vssd1
+ vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__o22a_1
XANTENNA__9255__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4571__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8697__B _3228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7855__A2 allocation.game.controller.drawBlock.state\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4746__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 allocation.game.lcdOutput.tft.remainingDelayTicks\[0\] vssd1 vssd1 vccd1 vccd1
+ net326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4841__A2 _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5730_ _1652_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5661_ _0769_ _0892_ _1585_ _1583_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__a31o_1
X_7400_ net251 net248 vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8380_ net148 _0471_ _0479_ vssd1 vssd1 vccd1 vccd1 _3841_ sky130_fd_sc_hd__and3_1
X_4612_ _0480_ _0542_ _0539_ net151 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoY\[7\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__9128__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5592_ _1513_ _1514_ _1516_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__and3_1
X_4543_ net106 vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__inv_2
X_7331_ allocation.game.cactus1size.lfsr1\[1\] allocation.game.cactus1size.lfsr2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7262_ allocation.game.controller.init_module.delay_counter\[1\] allocation.game.controller.init_module.delay_counter\[0\]
+ _2926_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6213_ _1042_ _1047_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__nor2_1
X_9001_ _4393_ _4394_ _4414_ _4449_ vssd1 vssd1 vccd1 vccd1 _4450_ sky130_fd_sc_hd__a31o_1
XANTENNA__9278__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4474_ net253 vssd1 vssd1 vccd1 vccd1 _4463_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7193_ allocation.game.dinoJump.count\[6\] allocation.game.dinoJump.count\[7\] vssd1
+ vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6144_ _2056_ _2068_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__nor2_1
X_6075_ net141 _0886_ net86 _0715_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__o22a_1
X_5026_ _0731_ _0949_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__or2_1
XANTENNA__6282__B2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6282__A1 _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6977_ allocation.game.scoreCounter.clock_div.counter\[17\] _2721_ net92 vssd1 vssd1
+ vccd1 vccd1 _2722_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_24_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5928_ _1852_ _1851_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__and2b_1
X_8716_ net164 net49 vssd1 vssd1 vccd1 vccd1 _4167_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5859_ _1735_ _1782_ _1783_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__nand3_1
X_8647_ _0635_ net142 _3602_ vssd1 vssd1 vccd1 vccd1 _4098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8731__B1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8578_ net47 _3256_ _4028_ _4026_ vssd1 vssd1 vccd1 vccd1 _4029_ sky130_fd_sc_hd__or4b_1
XANTENNA__5934__B _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7529_ _3054_ _3082_ _3138_ net246 vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4837__Y _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6491__A2_N _2234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6025__A1 _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6025__B2 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9092__RESET_B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5844__B _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6021__A _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5860__A _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8005__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7880_ allocation.game.controller.drawBlock.counter\[4\] _3415_ vssd1 vssd1 vccd1
+ vccd1 _3418_ sky130_fd_sc_hd__nand2_1
X_6900_ allocation.game.cactusDist.clock_div_inst0.counter\[1\] allocation.game.cactusDist.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__or2_1
X_6831_ allocation.game.cactus2size.clock_div_inst0.counter\[5\] allocation.game.cactus2size.clock_div_inst0.counter\[6\]
+ _2625_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6762_ net160 _2581_ _2582_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__nor3_1
X_8501_ _3949_ _3952_ _3278_ vssd1 vssd1 vccd1 vccd1 _3953_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9481_ clknet_leaf_7_clk _0388_ net193 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.v\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5713_ _0914_ _1637_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6693_ allocation.game.cactus1size.clock_div_inst1.counter\[1\] allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ allocation.game.cactus1size.clock_div_inst1.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2537_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5644_ _1519_ _1520_ _1511_ _1513_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__o211a_1
X_8432_ _3882_ _3884_ _3883_ vssd1 vssd1 vccd1 vccd1 _3885_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8411__A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8363_ _3574_ _3808_ _3823_ vssd1 vssd1 vccd1 vccd1 _3825_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7314_ allocation.game.controller.init_module.delay_counter\[19\] _2963_ net123 vssd1
+ vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5575_ _0831_ _1493_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout202_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8294_ net280 _3760_ vssd1 vssd1 vccd1 vccd1 _3761_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4526_ net234 _4455_ allocation.game.dinoJump.button vssd1 vssd1 vccd1 vccd1 _0464_
+ sky130_fd_sc_hd__and3_1
X_7245_ net264 allocation.game.dinoJump.next_dinoY\[5\] vssd1 vssd1 vccd1 vccd1 _2916_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7176_ _0472_ _2866_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6127_ _2049_ _2051_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout192_X net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _1981_ _1982_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__nor2_1
X_5009_ net60 _0932_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_29_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8305__B _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9443__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5049__A2 _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5360_ _0976_ _0989_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5291_ _1193_ _1213_ _1215_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7030_ _0446_ _2749_ _2752_ allocation.game.scoreCounter.bcd_tens\[1\] vssd1 vssd1
+ vccd1 vccd1 net24 sky130_fd_sc_hd__a31o_1
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4477__Y _0417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9316__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8981_ _0661_ net67 _4424_ _4429_ vssd1 vssd1 vccd1 vccd1 _4430_ sky130_fd_sc_hd__o211a_1
X_7932_ _0434_ _3453_ _3410_ vssd1 vssd1 vccd1 vccd1 _3455_ sky130_fd_sc_hd__o21a_1
XANTENNA__4653__B allocation.game.controller.drawBlock.y_end\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_7863_ allocation.game.controller.drawBlock.state\[3\] _2781_ _3402_ vssd1 vssd1
+ vccd1 vccd1 _3407_ sky130_fd_sc_hd__o21bai_1
XANTENNA__9466__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6814_ allocation.game.cactus2size.clock_div_inst0.counter\[7\] allocation.game.cactus2size.clock_div_inst0.counter\[6\]
+ allocation.game.cactus2size.clock_div_inst0.counter\[9\] allocation.game.cactus2size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__or4_1
X_7794_ net132 _3355_ vssd1 vssd1 vccd1 vccd1 _3356_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout152_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9533_ allocation.game.collides vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_6745_ allocation.game.cactus1size.clock_div_inst0.counter\[5\] _2569_ net154 vssd1
+ vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8141__A _0673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9464_ clknet_leaf_1_clk _0371_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6676_ _2523_ _2525_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_pixel\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8415_ net51 _3866_ vssd1 vssd1 vccd1 vccd1 _3868_ sky130_fd_sc_hd__or2_4
X_9395_ clknet_leaf_17_clk _0305_ net215 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5627_ net65 _1551_ _1549_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__a21o_1
X_8346_ _3807_ _3808_ vssd1 vssd1 vccd1 vccd1 _3809_ sky130_fd_sc_hd__and2b_1
X_5558_ _0787_ _1482_ _0786_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8277_ _3590_ _3742_ _3745_ net204 net429 vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__o32a_1
XFILLER_0_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4509_ net464 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7228_ net442 _2901_ _2903_ _0472_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__a211oi_1
X_5489_ _1411_ _1413_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7159_ allocation.game.lcdOutput.framebufferIndex\[12\] allocation.game.lcdOutput.framebufferIndex\[11\]
+ _2838_ _2859_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout65_A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5675__A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8456__A2 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9339__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9489__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5569__B _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4860_ _0782_ _0784_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__xnor2_1
X_4791_ _0565_ _0711_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6530_ _2428_ _2429_ _2415_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[8\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__5585__A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6461_ net218 _2378_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8200_ net105 _0691_ vssd1 vssd1 vccd1 vccd1 _3690_ sky130_fd_sc_hd__nand2_1
X_6392_ _2315_ vssd1 vssd1 vccd1 vccd1 allocation.game.collides sky130_fd_sc_hd__inv_2
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9180_ clknet_leaf_15_clk net338 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataShift\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5412_ _1334_ _1335_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__xor2_1
X_8131_ _0618_ _3630_ allocation.game.controller.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _3631_ sky130_fd_sc_hd__o21a_1
X_5343_ _1195_ _1212_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8062_ net231 _3562_ vssd1 vssd1 vccd1 vccd1 _3570_ sky130_fd_sc_hd__nand2_1
X_5274_ _0798_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__xnor2_2
X_7013_ allocation.game.bcd_ones\[1\] allocation.game.bcd_ones\[2\] allocation.game.bcd_ones\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7959__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8080__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8964_ _4000_ _4412_ _3998_ vssd1 vssd1 vccd1 vccd1 _4413_ sky130_fd_sc_hd__a21o_1
XANTENNA__7678__C net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7915_ allocation.game.controller.drawBlock.counter\[14\] _3439_ net95 vssd1 vssd1
+ vccd1 vccd1 _3443_ sky130_fd_sc_hd__o21ai_1
X_8895_ net262 _4255_ vssd1 vssd1 vccd1 vccd1 _4345_ sky130_fd_sc_hd__nand2_1
X_7846_ net426 _2975_ _3398_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__o21a_1
X_4989_ net78 _0904_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__or2_1
X_7777_ _3336_ _3338_ _3307_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5495__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9516_ net301 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_34_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6728_ allocation.game.cactus1size.clock_div_inst0.counter\[0\] _2557_ _2559_ allocation.game.cactus1size.clock_div_inst0.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__or4b_1
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9447_ clknet_leaf_11_clk _0397_ net201 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.drawDoneCactus
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6659_ net349 _2512_ _2514_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[31\]
+ sky130_fd_sc_hd__a21oi_1
X_9378_ clknet_leaf_9_clk _0288_ net196 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight2\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8329_ _3549_ _3778_ _3780_ vssd1 vssd1 vccd1 vccd1 _3793_ sky130_fd_sc_hd__nand3_1
XFILLER_0_30_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4880__A0 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout68_X net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_clk_X clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8601__A2 _3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5961_ _1840_ _1884_ _1885_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__nand3_1
X_4912_ _0830_ _0833_ _0836_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7700_ allocation.game.lcdOutput.framebufferIndex\[5\] net47 _3258_ vssd1 vssd1 vccd1
+ vccd1 _3262_ sky130_fd_sc_hd__a21o_1
X_8680_ net98 _4125_ _4130_ vssd1 vssd1 vccd1 vccd1 _4131_ sky130_fd_sc_hd__or3_1
X_5892_ _1814_ _1815_ _1813_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__a21bo_1
X_7631_ _0441_ _3189_ _3192_ vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__a21oi_2
X_4843_ _0758_ _0767_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__and2_4
XFILLER_0_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4774_ _0589_ _0595_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__xnor2_1
X_7562_ allocation.game.lcdOutput.tft.spi.counter\[2\] _2526_ vssd1 vssd1 vccd1 vccd1
+ _0250_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9301_ clknet_leaf_22_clk _0087_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6513_ _2417_ _2418_ net90 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7493_ _4463_ allocation.game.lcdOutput.tft.initSeqCounter\[4\] allocation.game.lcdOutput.tft.initSeqCounter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_9_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
X_6444_ _2334_ _2338_ _2366_ _2341_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__a31o_2
XFILLER_0_3_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9232_ clknet_leaf_22_clk _0029_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__7340__A2 _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout115_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7035__A _0417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6375_ allocation.game.cactusHeight1\[3\] _2279_ allocation.game.cactusHeight1\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__a21oi_1
X_9163_ clknet_leaf_15_clk _0225_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_9094_ clknet_leaf_14_clk _0190_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_8114_ _0643_ net164 _0654_ _0661_ vssd1 vssd1 vccd1 vccd1 _3615_ sky130_fd_sc_hd__o31ai_1
X_5326_ _1202_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8045_ _3518_ _0503_ vssd1 vssd1 vccd1 vccd1 _3554_ sky130_fd_sc_hd__nand2b_1
X_5257_ _0731_ _0947_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__xnor2_1
X_5188_ _1111_ _1112_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9034__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8947_ net97 _3694_ _4395_ net75 vssd1 vssd1 vccd1 vccd1 _4396_ sky130_fd_sc_hd__a22o_1
XANTENNA__8356__A1 _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8878_ _0467_ _3263_ _3811_ _4327_ vssd1 vssd1 vccd1 vccd1 _4328_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7829_ _2385_ _3384_ _3386_ _2360_ vssd1 vssd1 vccd1 vccd1 _3387_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5672__B net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout170 net174 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
Xfanout192 net200 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
Xfanout181 net188 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8044__B1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8595__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6024__A _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7554__S net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4490_ allocation.game.lcdOutput.tft.initSeqCounter\[2\] vssd1 vssd1 vccd1 vccd1
+ _0430_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6160_ _2082_ _2084_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5111_ _1022_ _1034_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__xnor2_1
X_6091_ _1978_ _2014_ _2013_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__a21o_1
X_5042_ _0964_ _0965_ _0937_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9057__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8586__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5103__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8801_ _3540_ _3760_ net261 vssd1 vssd1 vccd1 vccd1 _4251_ sky130_fd_sc_hd__a21oi_1
X_6993_ allocation.game.scoreCounter.clock_div.counter\[23\] _2730_ net92 vssd1 vssd1
+ vccd1 vccd1 _2732_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5944_ _1822_ _1865_ _1866_ _1868_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__a22o_1
X_8732_ net111 _0675_ _4180_ _4182_ vssd1 vssd1 vccd1 vccd1 _4183_ sky130_fd_sc_hd__o31ai_1
XANTENNA__8414__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4661__B allocation.game.controller.drawBlock.y_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8663_ _0669_ _4111_ _4113_ vssd1 vssd1 vccd1 vccd1 _4114_ sky130_fd_sc_hd__and3_1
X_5875_ _1798_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__and2b_1
X_4826_ _0750_ _0746_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__and2b_2
X_7614_ net232 allocation.game.game.score\[5\] net147 _2338_ vssd1 vssd1 vccd1 vccd1
+ _0278_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout232_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8594_ _4013_ _4027_ vssd1 vssd1 vccd1 vccd1 _4045_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7545_ _3149_ _3151_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4757_ allocation.game.controller.block_done net81 vssd1 vssd1 vccd1 vccd1 _0684_
+ sky130_fd_sc_hd__nor2_1
X_4688_ net225 _0613_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7849__B1 _3394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7476_ net364 net53 _3072_ _3091_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6427_ allocation.game.game.score\[1\] allocation.game.game.score\[0\] vssd1 vssd1
+ vccd1 vccd1 _2350_ sky130_fd_sc_hd__nor2_1
X_9215_ clknet_leaf_0_clk _0041_ net169 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9146_ clknet_leaf_9_clk _0210_ net196 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.x_dist\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6358_ allocation.game.cactusHeight1\[2\] _2278_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5309_ _0804_ _0833_ _0855_ _1018_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__a31o_1
X_9077_ clknet_leaf_14_clk _0173_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6289_ _2087_ _2200_ _2212_ _2213_ _2198_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__a2111o_1
X_8028_ net270 net163 _3526_ net241 net281 vssd1 vssd1 vccd1 vccd1 _3538_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4571__B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7068__B2 allocation.game.controller.drawBlock.y_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold4 allocation.game.lcdOutput.tft.spi.dataShift\[1\] vssd1 vssd1 vccd1 vccd1 net327
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9382__SET_B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6680__C _2526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5660_ _1538_ _1582_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4611_ _0540_ _0541_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8740__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5591_ _1490_ _1515_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4542_ _0471_ _0479_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nand2_1
X_7330_ allocation.game.cactusMove.drawDoneCactus _2974_ vssd1 vssd1 vccd1 vccd1 _2976_
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7261_ _2929_ _2930_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4473_ allocation.game.dinoJump.count\[20\] vssd1 vssd1 vccd1 vccd1 _4462_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6212_ _0797_ _1044_ _1048_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__a21oi_1
X_9000_ _4423_ _4439_ _4448_ vssd1 vssd1 vccd1 vccd1 _4449_ sky130_fd_sc_hd__and3_1
X_7192_ allocation.game.dinoJump.count\[6\] _2875_ allocation.game.dinoJump.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4937__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6143_ net110 _0900_ _2055_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4656__B allocation.game.controller.drawBlock.y_end\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6074_ _1985_ _1998_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__xor2_1
XANTENNA__7032__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _0731_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__nand2_1
XANTENNA__6282__A2 _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8559__B2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6976_ _2721_ net92 _2720_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_24_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5927_ _1849_ _1850_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__xnor2_1
X_8715_ net164 net49 vssd1 vssd1 vccd1 vccd1 _4166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5858_ _0777_ _0903_ _1733_ _1734_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8731__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout235_X net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8646_ _0685_ _2274_ vssd1 vssd1 vccd1 vccd1 _4097_ sky130_fd_sc_hd__nor2_1
X_4809_ _0558_ _0567_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__xnor2_4
X_5789_ net63 _1713_ _1712_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8577_ _4010_ _4016_ _4023_ _4027_ vssd1 vssd1 vccd1 vccd1 _4028_ sky130_fd_sc_hd__nand4_1
XFILLER_0_1_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7528_ net250 net252 _3050_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9222__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7459_ _3054_ _3073_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout95_A _3410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9129_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[23\] net185 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[23\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__7223__A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9372__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8798__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4566__B allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9510__295 vssd1 vssd1 vccd1 vccd1 _9510__295/HI net295 sky130_fd_sc_hd__conb_1
XANTENNA__4853__Y _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout50_X net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8722__B2 net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9408__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6021__B _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9061__RESET_B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4757__A allocation.game.controller.block_done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5860__B _0899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6830_ _2627_ _2628_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__nor2_1
XANTENNA__4923__C _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6761_ allocation.game.cactus1size.clock_div_inst0.counter\[11\] allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ _2578_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _1635_ _1636_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__xnor2_1
X_8500_ _4454_ _3939_ _0442_ _3313_ vssd1 vssd1 vccd1 vccd1 _3952_ sky130_fd_sc_hd__and4bb_1
X_9480_ clknet_leaf_7_clk _0387_ net195 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.v\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8713__A1 net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6692_ net153 _2530_ _2536_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_17_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5643_ _1567_ _1565_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__nand2b_1
X_8431_ net117 _3867_ vssd1 vssd1 vccd1 vccd1 _3884_ sky130_fd_sc_hd__nor2_1
XANTENNA__8411__B net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9245__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8362_ _3574_ _3808_ _3823_ vssd1 vssd1 vccd1 vccd1 _3824_ sky130_fd_sc_hd__nand3_1
X_5574_ _0801_ _0892_ _1498_ _1495_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7313_ net399 _2961_ _2964_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__o21a_1
X_4525_ net234 _4455_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8293_ net278 net275 vssd1 vssd1 vccd1 vccd1 _3760_ sky130_fd_sc_hd__or2_4
XFILLER_0_13_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7244_ net260 allocation.game.dinoJump.next_dinoY\[7\] vssd1 vssd1 vccd1 vccd1 _2915_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__9395__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7175_ allocation.game.dinoJump.count\[1\] _2864_ vssd1 vssd1 vccd1 vccd1 _2866_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6126_ _2032_ _2050_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_5_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6057_ _1940_ _1980_ _1979_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__a21oi_1
X_5008_ net60 _0932_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6959_ _2710_ net93 _2709_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__and3b_1
X_8629_ _4078_ _4079_ vssd1 vssd1 vccd1 vccd1 _4080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_10_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout98_X net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9118__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8943__A1 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9268__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5290_ _1157_ _1214_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8980_ _4428_ vssd1 vssd1 vccd1 vccd1 _4429_ sky130_fd_sc_hd__inv_2
X_7931_ allocation.game.controller.drawBlock.counter\[19\] _3409_ vssd1 vssd1 vccd1
+ vccd1 _3454_ sky130_fd_sc_hd__and2_1
X_7862_ allocation.game.controller.drawBlock.idx\[2\] _3402_ _3403_ _3406_ vssd1 vssd1
+ vccd1 vccd1 _0297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5748__A1 _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6813_ allocation.game.cactus2size.clock_div_inst0.counter\[1\] _2615_ allocation.game.cactus2size.clock_div_inst0.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__or3b_1
X_7793_ net130 net127 vssd1 vssd1 vccd1 vccd1 _3355_ sky130_fd_sc_hd__or2_1
X_9532_ net314 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
X_6744_ allocation.game.cactus1size.clock_div_inst0.counter\[5\] _2569_ vssd1 vssd1
+ vccd1 vccd1 _2571_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6675_ _2521_ _2524_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__nand2_1
X_9463_ clknet_leaf_18_clk _0370_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8414_ net50 _3866_ vssd1 vssd1 vccd1 vccd1 _3867_ sky130_fd_sc_hd__nand2_1
X_5626_ _1549_ _1550_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9394_ clknet_leaf_17_clk _0304_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8345_ _3547_ _3792_ _3806_ vssd1 vssd1 vccd1 vccd1 _3808_ sky130_fd_sc_hd__a21o_1
X_5557_ _0728_ _0778_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8276_ allocation.game.controller.state\[1\] _0437_ net240 _0436_ _3744_ vssd1 vssd1
+ vccd1 vccd1 _3745_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5488_ _1390_ _1409_ _1410_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__and3_1
X_4508_ net430 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
X_7227_ allocation.game.dinoJump.count\[16\] _2901_ vssd1 vssd1 vccd1 vccd1 _2903_
+ sky130_fd_sc_hd__nor2_1
X_7158_ _2848_ _2856_ _2858_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__a21oi_1
X_7089_ allocation.game.controller.drawBlock.x_start\[3\] _2772_ _2792_ allocation.game.controller.color\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__a22o_1
X_6109_ _1969_ _2006_ _2005_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__a21o_1
XANTENNA__9410__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5021__A _0938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8310__C1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8507__A _0401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7967__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9090__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7719__A2 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4790_ _0565_ _0711_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__xor2_4
XFILLER_0_28_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7557__S net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6460_ _2378_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5902__A1 _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6391_ _0462_ _2314_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5411_ _1335_ _1334_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__and2b_1
X_8130_ net223 _0617_ vssd1 vssd1 vccd1 vccd1 _3630_ sky130_fd_sc_hd__and2_1
X_5342_ _1246_ _1266_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8061_ net231 _3562_ vssd1 vssd1 vccd1 vccd1 _3569_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5273_ _0920_ _1196_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__and2_2
XFILLER_0_10_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7012_ allocation.game.bcd_ones\[0\] _2739_ _2744_ _2745_ vssd1 vssd1 vccd1 vccd1
+ net15 sky130_fd_sc_hd__o22a_1
XANTENNA__9433__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8963_ _4004_ _4411_ _4005_ vssd1 vssd1 vccd1 vccd1 _4412_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout262_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7914_ allocation.game.controller.drawBlock.counter\[14\] _3439_ vssd1 vssd1 vccd1
+ vccd1 _3442_ sky130_fd_sc_hd__and2_1
X_8894_ net36 _3811_ _4243_ _4216_ vssd1 vssd1 vccd1 vccd1 _4344_ sky130_fd_sc_hd__a31o_1
X_7845_ _3394_ _3397_ vssd1 vssd1 vccd1 vccd1 _3398_ sky130_fd_sc_hd__nand2_1
XANTENNA__4680__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8152__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4988_ _0903_ _0907_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__nor2_1
X_7776_ _3308_ _3334_ _3337_ vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__or3_1
X_9515_ net300 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_0_11_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6727_ allocation.game.cactus1size.clock_div_inst0.counter\[11\] allocation.game.cactus1size.clock_div_inst0.counter\[10\]
+ allocation.game.cactus1size.clock_div_inst0.counter\[13\] allocation.game.cactus1size.clock_div_inst0.counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__or4_1
X_9446_ clknet_leaf_9_clk _0396_ net195 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.drawDoneDino
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6658_ net349 _2512_ net146 vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9377_ clknet_leaf_9_clk _0287_ net196 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight2\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5609_ _1499_ _1500_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__xnor2_1
X_8328_ _3778_ _3780_ _3549_ vssd1 vssd1 vccd1 vccd1 _3792_ sky130_fd_sc_hd__a21o_1
X_6589_ allocation.game.cactusMove.count\[5\] _2468_ net149 vssd1 vssd1 vccd1 vccd1
+ _2471_ sky130_fd_sc_hd__o21ai_1
X_8259_ _2995_ _3731_ net54 vssd1 vssd1 vccd1 vccd1 _3732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8062__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9306__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4749__B net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5960_ _1836_ _1837_ _1839_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__a21o_1
X_4911_ _0834_ _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__nand2_1
X_5891_ _1813_ _1814_ _1815_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7630_ _0441_ net99 vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4842_ _0546_ _0571_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4773_ _0592_ _0696_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__or2_1
X_7561_ net360 net357 net256 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__mux2_1
X_9300_ clknet_leaf_22_clk _0086_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6512_ allocation.game.dinoJump.dinoDelay\[1\] allocation.game.dinoJump.dinoDelay\[0\]
+ allocation.game.dinoJump.dinoDelay\[2\] vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7492_ _4463_ net247 net249 _3052_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__or4_1
X_6443_ _2365_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__inv_2
X_9231_ clknet_leaf_0_clk _0028_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6374_ _4459_ _2292_ _2295_ net265 vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__o22a_1
X_9162_ clknet_leaf_15_clk _0224_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.data\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout108_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7035__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9093_ clknet_leaf_14_clk _0189_ net212 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_8113_ net142 _0644_ _0654_ _0661_ vssd1 vssd1 vccd1 vccd1 _3614_ sky130_fd_sc_hd__or4_1
X_5325_ _1016_ _1201_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__xor2_1
X_8044_ net107 _3552_ net244 vssd1 vssd1 vccd1 vccd1 _3553_ sky130_fd_sc_hd__o21a_1
X_5256_ _1179_ _1180_ _1178_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__o21ai_1
X_5187_ _1105_ _1109_ _1110_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__nor3_1
XANTENNA__4962__X _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8946_ _2312_ _2376_ vssd1 vssd1 vccd1 vccd1 _4395_ sky130_fd_sc_hd__or2_1
X_8877_ net266 _4308_ net41 vssd1 vssd1 vccd1 vccd1 _4327_ sky130_fd_sc_hd__a21o_1
XANTENNA__9329__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7828_ _2349_ _3385_ vssd1 vssd1 vccd1 vccd1 _3386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7759_ net68 net58 vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__nand2_4
XFILLER_0_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9479__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9429_ clknet_leaf_11_clk _0338_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout80_X net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 net184 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_4
Xfanout171 net174 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_4
Xfanout160 net162 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
XANTENNA__8044__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout193 net195 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8283__A1 allocation.game.controller.drawBlock.y_end\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7570__S _2526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5110_ _1022_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6090_ _1978_ _2013_ _2014_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5041_ _0937_ _0964_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8800_ net258 _4245_ vssd1 vssd1 vccd1 vccd1 _4250_ sky130_fd_sc_hd__xnor2_1
X_6992_ _2730_ _2731_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__nor2_1
X_8731_ net104 _4181_ net89 vssd1 vssd1 vccd1 vccd1 _4182_ sky130_fd_sc_hd__a21o_1
X_5943_ _1822_ _1865_ _1867_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5874_ _0728_ net103 _1027_ _1028_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__a2bb2o_1
X_8662_ net111 _4112_ _4107_ vssd1 vssd1 vccd1 vccd1 _4113_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4825_ _0710_ _0741_ _0748_ _0747_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__o31a_1
X_7613_ net232 allocation.game.game.score\[4\] net147 _2334_ vssd1 vssd1 vccd1 vccd1
+ _0277_ sky130_fd_sc_hd__a22o_1
X_8593_ net68 _3620_ _4039_ _4042_ vssd1 vssd1 vccd1 vccd1 _4044_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7544_ net253 _3039_ vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ net243 _0681_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__nand2_1
XANTENNA__5572__A2 _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4687_ net224 _0612_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__or2_1
X_7475_ _3020_ _3090_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6426_ _2348_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__inv_2
X_9214_ clknet_leaf_0_clk _0040_ net169 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6357_ net273 _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__nand2_1
X_9145_ clknet_leaf_18_clk net330 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_5308_ _1017_ _1026_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__xnor2_1
X_9076_ clknet_leaf_14_clk _0172_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6288_ allocation.game.controller.drawBlock.counter\[6\] _2195_ vssd1 vssd1 vccd1
+ vccd1 _2213_ sky130_fd_sc_hd__nor2_1
X_8027_ net270 net139 _3536_ net244 vssd1 vssd1 vccd1 vccd1 _3537_ sky130_fd_sc_hd__o211a_1
X_5239_ _1161_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_4_clk_X clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9151__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8929_ _4216_ _4244_ _4373_ net35 _4378_ vssd1 vssd1 vccd1 vccd1 _4379_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9515__300 vssd1 vssd1 vccd1 vccd1 _9515__300/HI net300 sky130_fd_sc_hd__conb_1
XFILLER_0_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5204__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 _0247_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload3_A clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output21_A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4610_ net258 allocation.game.controller.v\[7\] vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5590_ _1487_ _1489_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4541_ allocation.game.dinoJump.count\[9\] allocation.game.dinoJump.count\[11\] _0473_
+ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4472_ allocation.game.dinoJump.count\[18\] vssd1 vssd1 vccd1 vccd1 _4461_ sky130_fd_sc_hd__inv_2
X_7260_ net465 _2926_ net122 vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6211_ net63 _1058_ _1057_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__a21o_1
X_7191_ net419 _2875_ _2876_ _0472_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_42_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6142_ _0715_ net124 vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6073_ _1995_ _1997_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__xnor2_1
X_5024_ _0784_ _0947_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_0_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6975_ allocation.game.scoreCounter.clock_div.counter\[16\] allocation.game.scoreCounter.clock_div.counter\[15\]
+ _2717_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5926_ _0896_ _1744_ _1743_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__a21bo_1
X_8714_ net57 _3668_ _4163_ _4164_ vssd1 vssd1 vccd1 vccd1 _4165_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8645_ _4092_ _4095_ vssd1 vssd1 vccd1 vccd1 _4096_ sky130_fd_sc_hd__nand2_1
X_5857_ _1779_ _1781_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4808_ net80 _0731_ _0725_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__o21ai_1
X_8576_ _2517_ net51 vssd1 vssd1 vccd1 vccd1 _4027_ sky130_fd_sc_hd__xnor2_2
X_5788_ _1710_ _1711_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4739_ net220 allocation.game.cactusMove.x_dist\[7\] vssd1 vssd1 vccd1 vccd1 _0666_
+ sky130_fd_sc_hd__nor2_1
X_7527_ net248 _3074_ _3083_ _3119_ vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7458_ _3073_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6409_ allocation.game.game.score\[4\] _2330_ _2328_ vssd1 vssd1 vccd1 vccd1 _2332_
+ sky130_fd_sc_hd__o21a_1
X_7389_ net439 _2647_ _3014_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout88_A _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9128_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[22\] net185 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[22\] sky130_fd_sc_hd__dfrtp_1
X_9059_ clknet_leaf_20_clk allocation.game.dinoJump.next_dinoDelay\[5\] net192 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__4808__A1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7385__S _2973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5694__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8722__A2 _3228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7930__B1 _3409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9047__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4757__B net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9030__RESET_B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8961__A2 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6760_ allocation.game.cactus1size.clock_div_inst0.counter\[10\] _2578_ allocation.game.cactus1size.clock_div_inst0.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_18_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5711_ _0778_ net102 vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_18_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6691_ allocation.game.cactus1size.clock_div_inst1.counter\[1\] allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5642_ _1564_ _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__nand2_1
X_8430_ net114 _3868_ _3882_ _3880_ vssd1 vssd1 vccd1 vccd1 _3883_ sky130_fd_sc_hd__a31oi_2
X_8361_ allocation.game.controller.v\[6\] _0541_ _3562_ _3822_ vssd1 vssd1 vccd1 vccd1
+ _3823_ sky130_fd_sc_hd__o31a_1
X_5573_ _1495_ _1497_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__nor2_1
X_7312_ net123 _2963_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__nor2_1
X_4524_ net234 _4455_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__and2_2
X_8292_ net276 _3472_ vssd1 vssd1 vccd1 vccd1 _3759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7243_ _4462_ net144 _2912_ _2914_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__o31a_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7174_ net84 _2864_ _2865_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__and3_1
X_6125_ _2030_ _2031_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7330__Y _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6056_ _1940_ _1979_ _1980_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__and3_1
XANTENNA__7452__A2 _3066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5007_ _0858_ _0859_ _0861_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__o21ba_1
XANTENNA__4683__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6958_ allocation.game.scoreCounter.clock_div.counter\[10\] _2708_ vssd1 vssd1 vccd1
+ vccd1 _2710_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5909_ _1787_ _1832_ _1833_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__nand3_2
X_6889_ net437 _2665_ net152 vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__o21ai_1
X_8628_ _2520_ net57 vssd1 vssd1 vccd1 vccd1 _4079_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8559_ _4000_ _4002_ _4009_ net99 _4008_ vssd1 vssd1 vccd1 vccd1 _4010_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5689__A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6642__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7930_ net95 _3451_ _3453_ _3409_ allocation.game.controller.drawBlock.counter\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__a32o_1
X_7861_ _2781_ _3405_ _3400_ vssd1 vssd1 vccd1 vccd1 _3406_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4790__X _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9212__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6812_ allocation.game.cactus2size.clock_div_inst0.counter\[3\] allocation.game.cactus2size.clock_div_inst0.counter\[2\]
+ allocation.game.cactus2size.clock_div_inst0.counter\[5\] allocation.game.cactus2size.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__or4_1
XANTENNA__5748__A2 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7792_ _3287_ _3301_ _3310_ _3340_ _3353_ vssd1 vssd1 vccd1 vccd1 _3354_ sky130_fd_sc_hd__a311o_1
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6743_ _2569_ _2570_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__nor2_1
X_9531_ net313 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__9362__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6674_ net225 net223 net219 vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__and3_2
XFILLER_0_2_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9462_ clknet_leaf_18_clk _0369_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8413_ _3256_ _3863_ vssd1 vssd1 vccd1 vccd1 _3866_ sky130_fd_sc_hd__nor2_2
X_5625_ _1535_ _1547_ _1548_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__and3_1
X_9393_ clknet_leaf_17_clk _0303_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_8344_ _3547_ _3792_ _3806_ vssd1 vssd1 vccd1 vccd1 _3807_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5556_ _1430_ _1431_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__xnor2_1
X_8275_ net244 _3740_ _3743_ net163 net280 vssd1 vssd1 vccd1 vccd1 _3744_ sky130_fd_sc_hd__a32o_1
X_4507_ net432 vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
X_5487_ _1385_ _1403_ _1405_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7226_ allocation.game.dinoJump.count\[15\] _2900_ _2902_ vssd1 vssd1 vccd1 vccd1
+ _0165_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7157_ _2848_ _2849_ _2856_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__a21oi_1
X_7088_ allocation.game.controller.drawBlock.y_end\[3\] _2779_ _2803_ _2804_ vssd1
+ vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__a211o_1
X_6108_ _2004_ _2032_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6039_ _1861_ _1963_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8613__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4875__X _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9235__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9385__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6390_ _0617_ _2310_ _2312_ _2313_ _2277_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__a41o_1
X_5410_ _1284_ _1286_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5341_ _1248_ _1265_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__or2_1
X_8060_ net136 _3567_ _3566_ _3556_ vssd1 vssd1 vccd1 vccd1 _3568_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5272_ _0889_ _1196_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__and2_4
X_7011_ _0450_ allocation.game.bcd_ones\[3\] _2738_ vssd1 vssd1 vccd1 vccd1 _2745_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__4785__X _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8962_ net222 _3200_ _4409_ _4410_ vssd1 vssd1 vccd1 vccd1 _4411_ sky130_fd_sc_hd__o22a_1
X_7913_ net95 _3440_ _3441_ _3409_ allocation.game.controller.drawBlock.counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8893_ _4258_ _4342_ vssd1 vssd1 vccd1 vccd1 _4343_ sky130_fd_sc_hd__nor2_1
X_7844_ _2973_ _3393_ vssd1 vssd1 vccd1 vccd1 _3397_ sky130_fd_sc_hd__nor2_1
X_7775_ net51 net48 vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__nand2_1
X_9514_ net299 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
X_4987_ _0901_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__nand2_1
X_6726_ allocation.game.cactus1size.clock_div_inst0.counter\[7\] allocation.game.cactus1size.clock_div_inst0.counter\[6\]
+ allocation.game.cactus1size.clock_div_inst0.counter\[9\] allocation.game.cactus1size.clock_div_inst0.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9445_ clknet_leaf_11_clk _0354_ net202 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.cactusMovement
+ sky130_fd_sc_hd__dfrtp_1
X_6657_ _2512_ _2513_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[30\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6588_ allocation.game.cactusMove.count\[5\] _2468_ vssd1 vssd1 vccd1 vccd1 _2470_
+ sky130_fd_sc_hd__and2_1
XANTENNA__9108__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5608_ _1487_ _1532_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__and2_1
X_9376_ clknet_leaf_1_clk net325 net165 vssd1 vssd1 vccd1 vccd1 allocation.game.det
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8327_ _3789_ _3791_ allocation.game.controller.drawBlock.y_end\[4\] net201 vssd1
+ vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__o2bb2a_1
X_5539_ _1459_ _1462_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6400__B _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8258_ allocation.game.lcdOutput.tft.remainingDelayTicks\[18\] _2994_ vssd1 vssd1
+ vccd1 vccd1 _3731_ sky130_fd_sc_hd__nand2_1
XANTENNA__9258__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7209_ _0471_ _2888_ _2890_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__and3_1
X_8189_ _0691_ _3679_ net77 vssd1 vssd1 vccd1 vccd1 _3680_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8359__B1 allocation.game.controller.drawBlock.y_end\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5648__A1 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6309__Y _2234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4910_ _0831_ _0833_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _0712_ _0887_ _1768_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__a21o_1
X_4841_ _0760_ _0762_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_34_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7560_ net350 allocation.game.lcdOutput.tft.spi.data\[7\] net256 vssd1 vssd1 vccd1
+ vccd1 _0248_ sky130_fd_sc_hd__mux2_1
X_4772_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7491_ _3103_ _3104_ vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__xnor2_1
X_6511_ allocation.game.dinoJump.dinoDelay\[1\] allocation.game.dinoJump.dinoDelay\[0\]
+ allocation.game.dinoJump.dinoDelay\[2\] vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6442_ _2349_ _2364_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9230_ clknet_leaf_0_clk _0027_ net178 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_21_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9161_ clknet_leaf_19_clk _0223_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.tft_reset
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6373_ _2245_ _2296_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__and2_1
X_8112_ allocation.game.controller.drawBlock.x_end\[4\] net205 _3611_ _3613_ vssd1
+ vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9400__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9092_ clknet_leaf_14_clk _0188_ net215 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_5324_ _1016_ _1201_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__nand2_1
X_8043_ net265 net137 _3550_ _3551_ vssd1 vssd1 vccd1 vccd1 _3552_ sky130_fd_sc_hd__o22a_1
X_5255_ _1175_ _1177_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__xnor2_1
X_5186_ _1105_ _1109_ _1110_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__o21a_1
X_8945_ _2293_ _3275_ _4385_ vssd1 vssd1 vccd1 vccd1 _4394_ sky130_fd_sc_hd__a21o_1
X_8876_ _4313_ _4325_ vssd1 vssd1 vccd1 vccd1 _4326_ sky130_fd_sc_hd__nand2_1
XANTENNA__9002__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7827_ _2344_ _2357_ vssd1 vssd1 vccd1 vccd1 _3385_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7758_ _3293_ _3317_ _3318_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8610__B net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6709_ allocation.game.cactus1size.clock_div_inst1.counter\[7\] _2544_ allocation.game.cactus1size.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__a21oi_1
X_7689_ _3229_ _3250_ vssd1 vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__xor2_1
X_9428_ clknet_leaf_12_clk _0337_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9080__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9359_ clknet_leaf_12_clk _0008_ net204 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4866__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout172 net173 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_2
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4872__Y _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8073__A _4459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5697__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6321__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5040_ _0880_ _0882_ _0963_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6991_ allocation.game.scoreCounter.clock_div.counter\[22\] _2729_ net92 vssd1 vssd1
+ vccd1 vccd1 _2731_ sky130_fd_sc_hd__o21ai_1
X_5942_ _0741_ net102 _0908_ net103 vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__o22a_1
X_8730_ net111 _4180_ vssd1 vssd1 vccd1 vccd1 _4181_ sky130_fd_sc_hd__nor2_1
XANTENNA__5400__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8661_ _0673_ net98 _4104_ _4105_ vssd1 vssd1 vccd1 vccd1 _4112_ sky130_fd_sc_hd__o22a_1
X_5873_ _1796_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4824_ _0748_ _0709_ _0747_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_32_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8592_ _4032_ _4037_ _4039_ _4041_ vssd1 vssd1 vccd1 vccd1 _4043_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_28_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7612_ _4455_ allocation.game.game.score\[3\] net145 _2349_ vssd1 vssd1 vccd1 vccd1
+ _0276_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4755_ net243 _0681_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7543_ _3149_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout120_A _3181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7849__A2 _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4686_ net225 net221 vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__nor2_1
X_9213_ clknet_leaf_22_clk _0039_ net167 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_7474_ net253 allocation.game.lcdOutput.tft.initSeqCounter\[1\] _3021_ _3081_ _3089_
+ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__o311a_1
X_6425_ _2319_ _2346_ _2347_ _2330_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_45_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6356_ allocation.game.cactusHeight1\[3\] _2279_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__xnor2_4
X_9144_ clknet_leaf_18_clk _0208_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9075_ clknet_leaf_9_clk _0171_ net193 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoMovement
+ sky130_fd_sc_hd__dfrtp_2
X_5307_ _1183_ _1231_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__or2_1
X_8026_ _3534_ _3535_ net135 vssd1 vssd1 vccd1 vccd1 _3536_ sky130_fd_sc_hd__a21o_1
X_6287_ _2087_ _2200_ _2202_ allocation.game.controller.drawBlock.counter\[3\] _2211_
+ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__o221ai_1
X_5238_ _1160_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__and2_1
X_5169_ _1074_ _1091_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_3_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8928_ net35 _4373_ _4374_ _4377_ vssd1 vssd1 vccd1 vccd1 _4378_ sky130_fd_sc_hd__o22a_1
XANTENNA__9446__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8859_ net270 net43 vssd1 vssd1 vccd1 vccd1 _4309_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8670__C1 net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 allocation.game.lcdOutput.tft.remainingDelayTicks\[23\] vssd1 vssd1 vccd1 vccd1
+ net329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4540_ _0475_ _0476_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_10_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4471_ allocation.game.dinoJump.count\[8\] vssd1 vssd1 vccd1 vccd1 _4460_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6210_ _1063_ _2134_ _1061_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7190_ allocation.game.dinoJump.count\[6\] _2875_ vssd1 vssd1 vccd1 vccd1 _2876_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6141_ _2063_ _2064_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__xnor2_1
XANTENNA__9319__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6072_ _1957_ _1996_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__nand2_1
XANTENNA__4793__X _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5023_ _0784_ _0947_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6974_ allocation.game.scoreCounter.clock_div.counter\[15\] allocation.game.scoreCounter.clock_div.counter\[14\]
+ _2715_ allocation.game.scoreCounter.clock_div.counter\[16\] vssd1 vssd1 vccd1 vccd1
+ _2720_ sky130_fd_sc_hd__a31o_1
XANTENNA__5130__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8713_ net57 _3668_ _4149_ vssd1 vssd1 vccd1 vccd1 _4164_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5925_ _1765_ _1801_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5856_ _0769_ _0903_ _1779_ _1780_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_24_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8644_ _4093_ _4094_ vssd1 vssd1 vccd1 vccd1 _4095_ sky130_fd_sc_hd__nor2_1
X_4807_ net80 _0731_ _0725_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5787_ _1710_ _1711_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8575_ net229 net49 vssd1 vssd1 vccd1 vccd1 _4026_ sky130_fd_sc_hd__xor2_1
X_4738_ _0631_ _0639_ _0629_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7526_ net359 net53 _3129_ _3136_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4669_ _0596_ _0597_ _0586_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__a21o_1
X_7457_ _4463_ net251 vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6408_ allocation.game.game.score\[4\] _2330_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9127_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[21\] net185 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7388_ net282 net161 vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__nor2_2
X_6339_ _2254_ _2257_ _2262_ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_1_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_9058_ clknet_leaf_20_clk allocation.game.dinoJump.next_dinoDelay\[4\] net192 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[4\] sky130_fd_sc_hd__dfrtp_1
X_8009_ _0504_ _3518_ vssd1 vssd1 vccd1 vccd1 _3519_ sky130_fd_sc_hd__nand2_1
XANTENNA__4808__A2 _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8616__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout36_X net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8543__A_N net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7930__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5710_ net78 _0799_ _0908_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_18_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6690_ allocation.game.cactus1size.clock_div_inst1.counter\[0\] net153 _2534_ vssd1
+ vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__and3b_1
XFILLER_0_17_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5641_ _1517_ _1563_ _1562_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__o21ai_1
X_8360_ net231 _3562_ _3585_ vssd1 vssd1 vccd1 vccd1 _3822_ sky130_fd_sc_hd__o21ai_1
X_5572_ _0777_ _0885_ _1494_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__a21oi_1
X_7311_ allocation.game.controller.init_module.delay_counter\[18\] _2961_ vssd1 vssd1
+ vccd1 vccd1 _2963_ sky130_fd_sc_hd__and2_1
X_8291_ _0496_ _0524_ _3493_ _3756_ vssd1 vssd1 vccd1 vccd1 _3758_ sky130_fd_sc_hd__nand4_1
XANTENNA_clkbuf_leaf_3_clk_X clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4523_ _0454_ _0455_ _0460_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__nor3_1
X_7242_ net148 _0471_ _2911_ allocation.game.dinoJump.count\[20\] vssd1 vssd1 vccd1
+ vccd1 _2914_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9141__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7173_ allocation.game.dinoJump.count\[0\] net149 vssd1 vssd1 vccd1 vccd1 _2865_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6124_ _0761_ _0894_ _2028_ _2027_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__a31oi_2
XANTENNA__7988__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9291__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6055_ _1937_ _1939_ _1938_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__o21bai_1
X_5006_ _0854_ _0883_ _0930_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6957_ allocation.game.scoreCounter.clock_div.counter\[10\] _2708_ vssd1 vssd1 vccd1
+ vccd1 _2709_ sky130_fd_sc_hd__or2_1
XANTENNA__4970__Y _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5795__A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5908_ _1784_ _1786_ _1785_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__a21o_1
X_6888_ allocation.game.cactusDist.clock_div_inst1.counter\[12\] _2665_ vssd1 vssd1
+ vccd1 vccd1 _2666_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8627_ _2520_ net57 vssd1 vssd1 vccd1 vccd1 _4078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5839_ _1751_ _1756_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4726__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8558_ _4001_ _4002_ vssd1 vssd1 vccd1 vccd1 _4009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7509_ _3076_ _3119_ net245 vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8489_ _3890_ _3941_ _3896_ vssd1 vssd1 vccd1 vccd1 _3942_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9164__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7860_ allocation.game.controller.drawBlock.idx\[2\] _2761_ vssd1 vssd1 vccd1 vccd1
+ _3405_ sky130_fd_sc_hd__nor2_1
X_9528__322 vssd1 vssd1 vccd1 vccd1 net322 _9528__322/LO sky130_fd_sc_hd__conb_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6811_ allocation.game.cactus2size.clock_div_inst0.counter\[0\] allocation.game.cactus2size.clock_div_inst0.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__nand2_1
X_7791_ _3349_ _3352_ _3343_ vssd1 vssd1 vccd1 vccd1 _3353_ sky130_fd_sc_hd__o21a_1
XANTENNA__6504__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6742_ net435 _2567_ net154 vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__o21ai_1
X_9530_ net312 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
X_6673_ _2375_ _2521_ net219 vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__a21o_1
X_9461_ clknet_leaf_17_clk _0368_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9392_ clknet_leaf_17_clk _0302_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_8412_ _3864_ vssd1 vssd1 vccd1 vccd1 _3865_ sky130_fd_sc_hd__inv_2
X_5624_ _1535_ _1547_ _1548_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__a21oi_1
X_8343_ _3543_ _3571_ vssd1 vssd1 vccd1 vccd1 _3806_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9500__285 vssd1 vssd1 vccd1 vccd1 _9500__285/HI net285 sky130_fd_sc_hd__conb_1
X_5555_ _1478_ _1479_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout200_A allocation.game.cactus1size.clock_div_inst0.reset vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8274_ _0525_ net135 vssd1 vssd1 vccd1 vccd1 _3743_ sky130_fd_sc_hd__nand2_1
X_4506_ allocation.game.scoreCounter.bcd_tens\[0\] vssd1 vssd1 vccd1 vccd1 _0446_
+ sky130_fd_sc_hd__inv_2
X_5486_ _1390_ _1409_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__a21oi_1
X_7225_ _0472_ _2901_ vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__nor2_1
X_7156_ _0441_ _2857_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input5_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6107_ _2030_ _2031_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__or2_1
X_7087_ allocation.game.controller.drawBlock.x_end\[3\] _2777_ _2787_ allocation.game.controller.drawBlock.y_start\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__a22o_1
XANTENNA__9037__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6038_ _1816_ _1860_ _1859_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7989_ _3015_ net113 vssd1 vssd1 vccd1 vccd1 _3501_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_7_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8074__B1 _0541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8804__A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5340_ _1263_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__nand2_1
X_5271_ net79 _0891_ _0919_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__or3_1
X_7010_ allocation.game.bcd_ones\[0\] _2736_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__nor2_1
X_8961_ net224 net69 _4005_ _4073_ vssd1 vssd1 vccd1 vccd1 _4410_ sky130_fd_sc_hd__a211o_1
XANTENNA__8273__X _3742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7912_ _0433_ _3437_ vssd1 vssd1 vccd1 vccd1 _3441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8892_ _4249_ _4264_ _4335_ _4262_ vssd1 vssd1 vccd1 vccd1 _4342_ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4961__B _0706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7843_ allocation.game.cactusHeight2\[1\] _2976_ _3395_ vssd1 vssd1 vccd1 vccd1 _0288_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__4929__A1 _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4986_ _0903_ _0910_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout150_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7774_ net51 _3295_ _3335_ _3333_ vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__a31o_1
X_9513_ net298 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
X_6725_ allocation.game.cactus1size.clock_div_inst0.counter\[3\] allocation.game.cactus1size.clock_div_inst0.counter\[2\]
+ allocation.game.cactus1size.clock_div_inst0.counter\[5\] allocation.game.cactus1size.clock_div_inst0.counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9444_ clknet_leaf_11_clk _0353_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8977__A1_N net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6656_ net457 _2511_ net146 vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6587_ _2468_ _2469_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[4\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5607_ net82 _1486_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__or2_1
X_9375_ clknet_leaf_1_clk net324 net165 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.button
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8326_ net81 _2249_ _3785_ _3790_ vssd1 vssd1 vccd1 vccd1 _3791_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5538_ _1459_ _1462_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__and2b_1
X_8257_ net54 _3730_ _3027_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__o21ai_1
X_7208_ _2889_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__inv_2
X_5469_ _1197_ _1393_ _1392_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9102__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8188_ net112 _0658_ vssd1 vssd1 vccd1 vccd1 _3679_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7139_ net125 _2840_ allocation.game.lcdOutput.framebufferIndex\[15\] vssd1 vssd1
+ vccd1 vccd1 _2842_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5983__A _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4856__A0 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9352__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4840_ _0760_ _0763_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4771_ allocation.game.controller.drawBlock.y_start\[0\] allocation.game.controller.drawBlock.y_end\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__and2b_1
X_6510_ _0454_ _2414_ _2416_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[1\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__5584__A1 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7490_ _3042_ _3050_ _3053_ _3061_ vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6441_ _2363_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__inv_2
X_6372_ net259 _2292_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9160_ clknet_leaf_18_clk _0222_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8111_ allocation.game.controller.state\[7\] _3607_ _3612_ net243 vssd1 vssd1 vccd1
+ vccd1 _3613_ sky130_fd_sc_hd__a22o_1
X_5323_ _1246_ _1247_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__nand2_1
X_9091_ clknet_leaf_14_clk _0187_ net213 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8709__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8042_ _3530_ _3546_ net135 vssd1 vssd1 vccd1 vccd1 _3551_ sky130_fd_sc_hd__a21o_1
X_5254_ _0803_ _0842_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__nor2_1
X_5185_ _0969_ _0970_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout198_A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8589__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8944_ _2293_ _3276_ _4385_ _4392_ vssd1 vssd1 vccd1 vccd1 _4393_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8875_ _4458_ net128 _4324_ vssd1 vssd1 vccd1 vccd1 _4325_ sky130_fd_sc_hd__a21o_1
X_7826_ _2365_ _2371_ vssd1 vssd1 vccd1 vccd1 _3384_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9506__291 vssd1 vssd1 vccd1 vccd1 _9506__291/HI net291 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_35_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4969_ _0591_ _0697_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__and2_2
X_7757_ _3293_ _3318_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6708_ allocation.game.cactus1size.clock_div_inst1.counter\[7\] _2544_ _2546_ vssd1
+ vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7688_ allocation.game.lcdOutput.framebufferIndex\[5\] _3239_ net47 _3238_ vssd1
+ vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9427_ clknet_leaf_12_clk _0336_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_end\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_6639_ allocation.game.cactusMove.count\[24\] _2501_ vssd1 vssd1 vccd1 vccd1 _2502_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_22_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9225__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9358_ clknet_leaf_12_clk _0007_ net201 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_8309_ _4458_ net134 _3514_ _3774_ vssd1 vssd1 vccd1 vccd1 _3775_ sky130_fd_sc_hd__o211a_1
X_9289_ clknet_leaf_0_clk _0091_ net166 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__9375__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 _3461_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_4
Xfanout151 _0462_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout162 _2528_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
Xfanout195 net200 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net188 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
XANTENNA__8073__B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5697__B _0886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8752__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6321__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8268__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9338__283 vssd1 vssd1 vccd1 vccd1 _9338__283/HI net283 sky130_fd_sc_hd__conb_1
X_6990_ allocation.game.scoreCounter.clock_div.counter\[22\] _2729_ vssd1 vssd1 vccd1
+ vccd1 _2730_ sky130_fd_sc_hd__and2_1
XANTENNA__4792__A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5888__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _0762_ _0904_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__nor2_1
XANTENNA__8991__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8660_ _0675_ _4102_ _4106_ _4110_ vssd1 vssd1 vccd1 vccd1 _4111_ sky130_fd_sc_hd__a31o_1
X_5872_ _1745_ _1746_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4823_ _0716_ net110 vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8591_ _4041_ vssd1 vssd1 vccd1 vccd1 _4042_ sky130_fd_sc_hd__inv_2
X_7611_ net232 allocation.game.game.score\[2\] net146 _2356_ vssd1 vssd1 vccd1 vccd1
+ _0275_ sky130_fd_sc_hd__a22o_1
XANTENNA__9248__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4754_ _0663_ _0674_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7542_ net253 _3023_ _3037_ vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__and3_2
XFILLER_0_12_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7473_ _3041_ _3082_ _3088_ _3087_ allocation.game.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__a311o_1
X_4685_ net230 _0612_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__or2_1
X_9212_ clknet_leaf_0_clk _0034_ net175 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst1.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6424_ allocation.game.game.score\[3\] _2329_ _2328_ vssd1 vssd1 vccd1 vccd1 _2347_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__9398__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6355_ allocation.game.cactusHeight1\[1\] allocation.game.cactusHeight1\[0\] allocation.game.cactusHeight1\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__a21o_2
XANTENNA__4967__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9143_ clknet_leaf_18_clk _0207_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_5306_ _1027_ _1182_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__and2_1
X_9074_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[20\] net190 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6286_ allocation.game.controller.drawBlock.counter\[3\] _2202_ _2204_ allocation.game.controller.drawBlock.counter\[2\]
+ _2210_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_12_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8025_ _3530_ _3533_ vssd1 vssd1 vccd1 vccd1 _3535_ sky130_fd_sc_hd__or2_1
X_5237_ _1150_ _1157_ _1159_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5168_ _0853_ _1092_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__or2_1
X_5099_ _0772_ _0750_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5798__A _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8927_ net41 _3542_ _4375_ _3523_ _4376_ vssd1 vssd1 vccd1 vccd1 _4377_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8858_ net270 net43 vssd1 vssd1 vccd1 vccd1 _4308_ sky130_fd_sc_hd__nor2_1
X_7809_ net96 _3321_ _3370_ vssd1 vssd1 vccd1 vccd1 _3371_ sky130_fd_sc_hd__o21ai_1
X_8789_ net40 _4220_ vssd1 vssd1 vccd1 vccd1 _4239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8349__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7 _0209_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8084__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__8812__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4470_ net262 vssd1 vssd1 vccd1 vccd1 _4459_ sky130_fd_sc_hd__inv_2
XANTENNA__7700__A2 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6140_ _2063_ _2064_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6071_ _1954_ _1956_ _1955_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5022_ net80 _0782_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_0_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6973_ net424 _2717_ _2719_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9070__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5924_ _1843_ _1847_ _1811_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__o21a_1
X_8712_ _3208_ _3672_ _4159_ _4162_ vssd1 vssd1 vccd1 vccd1 _4163_ sky130_fd_sc_hd__a211o_1
X_5855_ net87 _0907_ _1778_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_24_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8643_ net257 _3248_ vssd1 vssd1 vccd1 vccd1 _4094_ sky130_fd_sc_hd__and2_1
X_4806_ _0724_ net72 vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5786_ _1651_ _1657_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8574_ _4010_ _4024_ _4006_ vssd1 vssd1 vccd1 vccd1 _4025_ sky130_fd_sc_hd__a21oi_1
X_7525_ _3133_ _3135_ net53 vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4737_ net220 allocation.game.cactusMove.x_dist\[7\] vssd1 vssd1 vccd1 vccd1 _0664_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_47_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4668_ _0586_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__nand2b_2
X_7456_ net368 _0233_ _3065_ _3072_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout116_X net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6407_ allocation.game.game.score\[3\] _2329_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4599_ _0502_ _0531_ net106 vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__a21oi_1
X_9126_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[20\] net185 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[20\] sky130_fd_sc_hd__dfrtp_1
X_7387_ allocation.game.cactusMove.x_dist\[7\] _2976_ _3013_ vssd1 vssd1 vccd1 vccd1
+ _0215_ sky130_fd_sc_hd__a21bo_1
X_6338_ net272 _2253_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__nand2_1
X_6269_ _2066_ _2078_ _2097_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__and3_1
X_9057_ clknet_leaf_2_clk allocation.game.dinoJump.next_dinoDelay\[3\] net191 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[3\] sky130_fd_sc_hd__dfrtp_1
X_8008_ _3504_ _3507_ _3517_ vssd1 vssd1 vccd1 vccd1 _3518_ sky130_fd_sc_hd__or3_1
XANTENNA__9413__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5991__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9093__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7382__B1 _2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _1553_ _1558_ _1560_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__a21bo_1
X_5571_ net71 _0892_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7310_ net417 _2959_ _2962_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__o21a_1
X_8290_ _0496_ _0524_ _3493_ _3756_ vssd1 vssd1 vccd1 vccd1 _3757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4522_ _0456_ _0457_ _0458_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7241_ net455 net144 _2912_ _2913_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__a22o_1
X_7172_ allocation.game.dinoJump.count\[0\] net149 vssd1 vssd1 vccd1 vccd1 _2864_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9436__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6123_ _2038_ _2046_ _2047_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__and3_1
XANTENNA_clkload15_A clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6054_ _1975_ _1978_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__nand2_1
X_5005_ _0884_ _0929_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__nor2_1
XANTENNA__4964__B _0886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5141__A _0754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8937__A1 _0401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9275__SET_B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6956_ _2392_ _2704_ _2707_ net479 net93 vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5907_ _1828_ _1831_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6887_ net159 _2664_ _2665_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5838_ _1762_ _1761_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8626_ net217 _2524_ _4030_ _4052_ _4076_ vssd1 vssd1 vccd1 vccd1 _4077_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8557_ net74 _4007_ vssd1 vssd1 vccd1 vccd1 _4008_ sky130_fd_sc_hd__nand2_1
X_5769_ _1689_ _1691_ _1693_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7508_ _3076_ _3119_ vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8488_ _3321_ _3325_ _3867_ vssd1 vssd1 vccd1 vccd1 _3941_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7439_ net251 _3045_ net248 vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9109_ clknet_leaf_6_clk allocation.game.cactusMove.n_count\[3\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6313__C _0673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9309__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9459__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8919__A1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8919__B2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6810_ net402 net161 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7790_ _3333_ _3351_ _3336_ vssd1 vssd1 vccd1 vccd1 _3352_ sky130_fd_sc_hd__a21boi_1
XANTENNA__6504__B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6741_ allocation.game.cactus1size.clock_div_inst0.counter\[3\] allocation.game.cactus1size.clock_div_inst0.counter\[4\]
+ _2566_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6672_ _2375_ _2521_ _2522_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_pixel\[6\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9460_ clknet_leaf_17_clk _0367_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6158__A1 _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9391_ clknet_leaf_17_clk _0301_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_8411_ net47 net46 vssd1 vssd1 vccd1 vccd1 _3864_ sky130_fd_sc_hd__or2_2
X_5623_ _1502_ _1503_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__xnor2_1
X_8342_ _3798_ _3805_ allocation.game.controller.drawBlock.y_end\[5\] net201 vssd1
+ vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5554_ _1473_ _1476_ _1477_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9535__316 vssd1 vssd1 vccd1 vccd1 _9535__316/HI net316 sky130_fd_sc_hd__conb_1
XFILLER_0_48_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8273_ net107 _3741_ net241 vssd1 vssd1 vccd1 vccd1 _3742_ sky130_fd_sc_hd__o21a_1
X_4505_ allocation.game.scoreCounter.bcd_tens\[1\] vssd1 vssd1 vccd1 vccd1 _0445_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5485_ _1343_ _1362_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__xnor2_1
X_7224_ allocation.game.dinoJump.count\[15\] _2900_ vssd1 vssd1 vccd1 vccd1 _2901_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4975__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7155_ allocation.game.lcdOutput.framebufferIndex\[10\] allocation.game.lcdOutput.framebufferIndex\[9\]
+ _2834_ _2838_ _2855_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__a32o_1
XANTENNA__8083__A1 allocation.game.controller.drawBlock.y_start\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6106_ _1999_ _2001_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__xnor2_1
X_7086_ allocation.game.controller.color\[11\] _2786_ vssd1 vssd1 vccd1 vccd1 _2803_
+ sky130_fd_sc_hd__and2_1
X_6037_ _1945_ _1961_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7988_ net244 _3497_ _3498_ _3499_ vssd1 vssd1 vccd1 vccd1 _3500_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6939_ allocation.game.scoreCounter.clock_div.counter\[0\] allocation.game.scoreCounter.clock_div.counter\[1\]
+ allocation.game.scoreCounter.clock_div.counter\[2\] vssd1 vssd1 vccd1 vccd1 _2699_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8609_ _4054_ _4055_ _4057_ _4059_ _4056_ vssd1 vssd1 vccd1 vccd1 _4060_ sky130_fd_sc_hd__o41a_1
XFILLER_0_49_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4580__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8310__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout96_X net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9049__RESET_B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_X clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7585__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9131__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9281__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5270_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7171__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4795__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8960_ net224 net69 _4056_ _4059_ vssd1 vssd1 vccd1 vccd1 _4409_ sky130_fd_sc_hd__o211a_1
X_7911_ _3439_ vssd1 vssd1 vccd1 vccd1 _3440_ sky130_fd_sc_hd__inv_2
X_8891_ _3294_ _3871_ _4332_ _4340_ _3931_ vssd1 vssd1 vccd1 vccd1 _4341_ sky130_fd_sc_hd__a32o_1
XANTENNA__6379__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7842_ _0437_ _2975_ _3396_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__o21ai_1
X_4985_ net102 _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__nor2_1
XANTENNA__5051__A1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7773_ _3334_ vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__inv_2
X_9512_ net297 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XANTENNA_fanout143_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6724_ net339 _2554_ _2556_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__a21oi_1
X_9443_ clknet_leaf_11_clk _0352_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6655_ allocation.game.cactusMove.count\[30\] _2511_ vssd1 vssd1 vccd1 vccd1 _2512_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6586_ net481 _2466_ net149 vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_30_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5606_ _1529_ _1530_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__and2b_1
X_9374_ clknet_leaf_1_clk net3 net165 vssd1 vssd1 vccd1 vccd1 allocation.game.sync0
+ sky130_fd_sc_hd__dfrtp_1
X_8325_ _2300_ net100 _2411_ _3523_ _3633_ vssd1 vssd1 vccd1 vccd1 _3790_ sky130_fd_sc_hd__o221a_1
X_5537_ _1434_ _1460_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8256_ allocation.game.lcdOutput.tft.remainingDelayTicks\[16\] _2993_ vssd1 vssd1
+ vccd1 vccd1 _3730_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7207_ allocation.game.dinoJump.count\[9\] allocation.game.dinoJump.count\[10\] _2885_
+ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__and3_1
X_5468_ _0846_ _1198_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__xnor2_1
X_8187_ net431 net207 _3678_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__o21ba_1
X_5399_ _1320_ _1322_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__xnor2_1
X_7138_ net125 _2840_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__nand2_1
X_7069_ _2756_ _2768_ _2780_ _2788_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__o22a_1
XANTENNA__9154__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout56_A net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5983__B _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5281__A1 _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9419__Q allocation.game.controller.drawBlock.y_start\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4770_ _0695_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7166__A _0401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6440_ _2353_ _2356_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__nor2_1
XANTENNA__4544__B1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9027__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6371_ _2292_ _2294_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__nor2_1
X_5322_ _1242_ _1245_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__or2_1
X_8110_ _0687_ _2274_ vssd1 vssd1 vccd1 vccd1 _3612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9090_ clknet_leaf_14_clk _0186_ net215 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.init_module.delay_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8041_ _3530_ _3549_ vssd1 vssd1 vccd1 vccd1 _3550_ sky130_fd_sc_hd__nor2_1
X_5253_ _1175_ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__or2_1
X_5184_ _1106_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__and2_1
X_8943_ net44 _4390_ _4391_ vssd1 vssd1 vccd1 vccd1 _4392_ sky130_fd_sc_hd__a21oi_1
X_8874_ _4314_ _4315_ _4323_ vssd1 vssd1 vccd1 vccd1 _4324_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7825_ net234 allocation.game.bcd_ones\[3\] vssd1 vssd1 vccd1 vccd1 _3383_ sky130_fd_sc_hd__or2_1
XANTENNA__7628__X _3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4968_ _0798_ _0889_ net86 vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__nor3_4
XFILLER_0_4_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7756_ net50 net48 vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__or2_2
XFILLER_0_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4899_ net82 _0822_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6707_ allocation.game.cactus1size.clock_div_inst1.counter\[7\] _2544_ net159 vssd1
+ vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7687_ net47 vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9426_ clknet_leaf_8_clk _0335_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_start\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6638_ _2501_ net150 _2500_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[23\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_22_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9357_ clknet_leaf_11_clk _0006_ net202 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_8308_ _3504_ _3513_ net134 vssd1 vssd1 vccd1 vccd1 _3774_ sky130_fd_sc_hd__o21ai_1
X_6569_ allocation.game.cactusMove.count\[21\] allocation.game.cactusMove.count\[20\]
+ allocation.game.cactusMove.count\[23\] allocation.game.cactusMove.count\[22\] vssd1
+ vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__or4_1
XANTENNA__7804__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9288_ clknet_leaf_1_clk _0103_ net166 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_8239_ allocation.game.lcdOutput.tft.remainingDelayTicks\[10\] _2989_ vssd1 vssd1
+ vccd1 vccd1 _3719_ sky130_fd_sc_hd__xor2_1
XANTENNA__8029__A1 allocation.game.controller.drawBlock.y_start\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xfanout163 _2412_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_4
Xfanout174 net200 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
Xfanout141 _0713_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout152 net157 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
Xfanout196 net198 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_4
Xfanout185 net187 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4882__B _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9064__RESET_B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7228__C1 _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7243__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4792__B _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5888__B _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5940_ _0741_ _0908_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7610_ _4455_ allocation.game.game.score\[1\] net145 _2353_ vssd1 vssd1 vccd1 vccd1
+ _0274_ sky130_fd_sc_hd__o22a_1
X_5871_ _1766_ _1777_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__a21bo_1
X_4822_ _0715_ _0724_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8590_ net75 _4038_ _4040_ _4032_ vssd1 vssd1 vccd1 vccd1 _4041_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4753_ _0663_ net105 vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7541_ net254 _3148_ _3147_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7472_ net249 _3052_ _3083_ net246 vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__o211a_1
X_4684_ net227 net226 vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__or2_2
X_6423_ _2325_ _2345_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__or2_1
X_9211_ _0149_ _0408_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6354_ allocation.game.cactusHeight1\[1\] allocation.game.cactusHeight1\[0\] vssd1
+ vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__nand2_2
X_9142_ clknet_leaf_18_clk _0206_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_5305_ _1229_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__inv_2
X_9073_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[19\] net189 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[19\] sky130_fd_sc_hd__dfrtp_1
X_6285_ allocation.game.controller.drawBlock.counter\[2\] _2204_ _2205_ _2206_ _2209_
+ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__o2111ai_1
X_8024_ _3530_ _3533_ vssd1 vssd1 vccd1 vccd1 _3534_ sky130_fd_sc_hd__nand2_1
X_5236_ _0924_ _1155_ _1153_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ _0829_ _0852_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__nor2_1
X_5098_ _0750_ _0772_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__and2b_1
XANTENNA__5798__B net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8926_ _3523_ _4375_ net44 vssd1 vssd1 vccd1 vccd1 _4376_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_9_Left_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8195__B1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8857_ net266 net40 vssd1 vssd1 vccd1 vccd1 _4307_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7808_ net96 net74 vssd1 vssd1 vccd1 vccd1 _3370_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8788_ _4222_ _4236_ _4237_ vssd1 vssd1 vccd1 vccd1 _4238_ sky130_fd_sc_hd__o21a_1
X_7739_ _3291_ _3295_ _3297_ _3290_ vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__o31a_1
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9342__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9409_ clknet_leaf_17_clk _0319_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5054__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8365__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 allocation.game.lcdOutput.tft.spi.dataShift\[7\] vssd1 vssd1 vccd1 vccd1 net331
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8973__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9522__307 vssd1 vssd1 vccd1 vccd1 _9522__307/HI net307 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_26_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7709__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6070_ _1951_ _1990_ _1991_ _1993_ _1994_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__a32o_1
XANTENNA__8661__A1 _0673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5021_ _0938_ _0945_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9215__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6972_ allocation.game.scoreCounter.clock_div.counter\[15\] _2717_ net92 vssd1 vssd1
+ vccd1 vccd1 _2719_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8711_ _4160_ _4161_ vssd1 vssd1 vccd1 vccd1 _4162_ sky130_fd_sc_hd__nand2_1
X_5923_ _1811_ _1847_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__xor2_1
X_5854_ net87 _0907_ _1778_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__nand3_1
XANTENNA__9365__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8642_ net257 net47 vssd1 vssd1 vccd1 vccd1 _4093_ sky130_fd_sc_hd__nor2_1
X_8573_ _4015_ _4020_ _4021_ _4022_ vssd1 vssd1 vccd1 vccd1 _4024_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4805_ _0729_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5785_ _1702_ _1707_ _1708_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7524_ net246 _3101_ _3134_ _3102_ _3060_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__a32o_1
X_4736_ _0651_ _0652_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4667_ allocation.game.controller.drawBlock.y_end\[3\] allocation.game.controller.drawBlock.y_start\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7455_ _3067_ _3068_ _3071_ net53 vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__o211ai_2
X_6406_ allocation.game.game.score\[2\] allocation.game.game.score\[1\] allocation.game.game.score\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__and3_1
X_7386_ allocation.game.cactusMove.x_dist\[6\] _2975_ _3013_ vssd1 vssd1 vccd1 vccd1
+ _0214_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout109_X net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4598_ _0491_ _0492_ _0501_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__nand3_1
X_6337_ net278 _2260_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__and2_1
X_9125_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[19\] net184 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[19\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__8101__B1 _2516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6268_ _2101_ _2192_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__nand2_1
X_9056_ clknet_leaf_2_clk allocation.game.dinoJump.next_dinoDelay\[2\] net191 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[2\] sky130_fd_sc_hd__dfrtp_1
X_8007_ _4458_ allocation.game.controller.v\[3\] vssd1 vssd1 vccd1 vccd1 _3517_ sky130_fd_sc_hd__nor2_1
X_5219_ _1124_ _1142_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__or2_1
X_6199_ _1424_ _2123_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__and2_1
X_8909_ _4357_ _4320_ vssd1 vssd1 vccd1 vccd1 _4359_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7915__B1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_22_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4660__A_N allocation.game.controller.drawBlock.y_start\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9238__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9388__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6343__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7906__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7382__A1 _3008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5570_ _0777_ _0885_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4521_ allocation.game.dinoJump.dinoDelay\[14\] allocation.game.dinoJump.dinoDelay\[17\]
+ allocation.game.dinoJump.dinoDelay\[16\] allocation.game.dinoJump.dinoDelay\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__or4b_1
X_7240_ allocation.game.dinoJump.count\[19\] _2909_ vssd1 vssd1 vccd1 vccd1 _2913_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7171_ net144 _0519_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6122_ _2035_ _2037_ _2036_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__a21o_1
XANTENNA__7621__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6053_ _1975_ _1976_ _1977_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__nand3_1
X_5004_ _0924_ _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4964__C _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8398__B1 allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8733__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6955_ _2392_ _2704_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5906_ _1828_ _1829_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6886_ allocation.game.cactusDist.clock_div_inst1.counter\[11\] allocation.game.cactusDist.clock_div_inst1.counter\[10\]
+ _2661_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__and3_1
X_8625_ _4067_ _4075_ _4071_ _4060_ vssd1 vssd1 vccd1 vccd1 _4076_ sky130_fd_sc_hd__o2bb2a_1
X_5837_ net63 _1713_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__xnor2_1
X_8556_ _0614_ _2374_ _3674_ net221 vssd1 vssd1 vccd1 vccd1 _4007_ sky130_fd_sc_hd__a22o_1
X_5768_ _0901_ _1642_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__xnor2_1
X_4719_ net228 _0644_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__nand2_1
X_8487_ _3362_ _3939_ vssd1 vssd1 vccd1 vccd1 _3940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7507_ net253 _3041_ net250 vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__a21oi_2
X_5699_ net88 _0892_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__nand2_1
X_7438_ _4463_ _3053_ _3051_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7369_ net376 _2995_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9108_ clknet_leaf_6_clk allocation.game.cactusMove.n_count\[2\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout86_A _0891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9039_ clknet_leaf_7_clk _0164_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8627__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8643__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout41_X net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9060__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8818__A net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6338__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8553__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5602__A1 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6740_ _2567_ _2568_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6671_ net225 _2521_ net221 vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9390_ clknet_leaf_17_clk _0300_ net208 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8410_ net49 net47 vssd1 vssd1 vccd1 vccd1 _3863_ sky130_fd_sc_hd__or2_1
X_5622_ _1545_ _1546_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8341_ net81 _2243_ _3803_ _3804_ vssd1 vssd1 vccd1 vccd1 _3805_ sky130_fd_sc_hd__o211a_1
X_5553_ _1473_ _1476_ _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4504_ allocation.game.controller.drawBlock.idx\[1\] vssd1 vssd1 vccd1 vccd1 _0444_
+ sky130_fd_sc_hd__inv_2
XANTENNA__9403__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8272_ _0525_ net137 _3740_ vssd1 vssd1 vccd1 vccd1 _3741_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5484_ _1406_ _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__nand2_1
X_7223_ net150 _2882_ _2899_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7154_ _2838_ _2855_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6105_ _1858_ _2029_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__nand2_1
X_7085_ _2794_ _2797_ vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__nand2b_1
X_6036_ _1958_ _1959_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__xnor2_1
X_7987_ allocation.game.collision.dinoY\[2\] net163 _3491_ net241 vssd1 vssd1 vccd1
+ vccd1 _3499_ sky130_fd_sc_hd__a22o_1
X_6938_ allocation.game.scoreCounter.clock_div.counter\[0\] net381 _2698_ vssd1 vssd1
+ vccd1 vccd1 _0116_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6869_ allocation.game.cactusDist.clock_div_inst1.counter\[4\] _2651_ allocation.game.cactusDist.clock_div_inst1.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8608_ net229 _3237_ _4058_ vssd1 vssd1 vccd1 vccd1 _4059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9083__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8539_ allocation.game.lcdOutput.framebufferIndex\[0\] _3285_ _3357_ _3278_ vssd1
+ vssd1 vccd1 vccd1 _3991_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_38_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4580__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout89_X net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8782__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5899__A1 _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6068__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7910_ _0433_ _3437_ vssd1 vssd1 vccd1 vccd1 _3439_ sky130_fd_sc_hd__nor2_1
X_8890_ net119 net66 _3292_ _3875_ vssd1 vssd1 vccd1 vccd1 _4340_ sky130_fd_sc_hd__a31o_1
X_7841_ _3393_ _3395_ vssd1 vssd1 vccd1 vccd1 _3396_ sky130_fd_sc_hd__nand2_1
X_4984_ net78 _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__or2_1
X_7772_ _3317_ _3325_ vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9511_ net296 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_6723_ net339 _2554_ net152 vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9442_ clknet_leaf_15_clk _0351_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_6654_ _2511_ net150 _2510_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[29\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5605_ _1527_ _1528_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__or2_1
XANTENNA__5147__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6585_ allocation.game.cactusMove.count\[3\] allocation.game.cactusMove.count\[4\]
+ _2465_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__and3_1
X_9373_ clknet_leaf_14_clk _0004_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8324_ _3479_ _3788_ allocation.game.controller.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _3789_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5536_ _1434_ _1460_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__and2_1
X_5467_ _0846_ _1198_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__nand2_1
X_8255_ _3727_ _3729_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__or2_1
X_7206_ allocation.game.dinoJump.count\[10\] _2886_ vssd1 vssd1 vccd1 vccd1 _2888_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_44_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8186_ _0660_ net77 _3672_ _0683_ _3677_ vssd1 vssd1 vccd1 vccd1 _3678_ sky130_fd_sc_hd__o221a_1
X_5398_ _1322_ _1320_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__nand2b_1
X_7137_ allocation.game.lcdOutput.framebufferIndex\[12\] allocation.game.lcdOutput.framebufferIndex\[13\]
+ _2839_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__and3_1
X_7068_ allocation.game.controller.color\[8\] _2786_ _2787_ allocation.game.controller.drawBlock.y_start\[0\]
+ _2784_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__a221o_1
XANTENNA__4992__Y _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6019_ _1927_ _1928_ _1907_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8368__A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7191__C1 _0472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4544__A1 _4459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6370_ allocation.game.cactusHeight1\[5\] _2291_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5321_ _1242_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8040_ _3547_ _3548_ vssd1 vssd1 vccd1 vccd1 _3549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5252_ _1134_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5183_ _1105_ _1107_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8942_ net44 _4390_ _2300_ vssd1 vssd1 vccd1 vccd1 _4391_ sky130_fd_sc_hd__o21a_1
X_8873_ _4317_ _4322_ _4316_ vssd1 vssd1 vccd1 vccd1 _4323_ sky130_fd_sc_hd__a21o_1
X_7824_ allocation.game.bcd_ones\[2\] _2369_ _3382_ net146 vssd1 vssd1 vccd1 vccd1
+ _0283_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4967_ net86 vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__inv_2
X_7755_ net68 net56 vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4898_ net82 _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__and2_1
X_7686_ _3244_ _3246_ _3242_ vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__o21ai_2
X_6706_ _2544_ _2545_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__nor2_1
X_9425_ clknet_leaf_12_clk _0334_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_start\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_6637_ allocation.game.cactusMove.count\[23\] allocation.game.cactusMove.count\[22\]
+ _2497_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9356_ clknet_leaf_12_clk _0005_ net206 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_6568_ allocation.game.cactusMove.count\[12\] allocation.game.cactusMove.count\[14\]
+ allocation.game.cactusMove.count\[15\] allocation.game.cactusMove.count\[13\] vssd1
+ vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__or4bb_1
X_8307_ _3769_ _3771_ _3772_ net241 vssd1 vssd1 vccd1 vccd1 _3773_ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5519_ _1196_ _1443_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__nand2_1
XANTENNA__7804__B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8277__A2 _3742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6499_ _0419_ _0681_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9287_ clknet_leaf_1_clk _0102_ net165 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_1_clk_X clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9121__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8238_ _2989_ _3717_ _3718_ net55 vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__a22oi_1
X_8169_ _3662_ vssd1 vssd1 vccd1 vccd1 _3663_ sky130_fd_sc_hd__inv_2
Xfanout131 allocation.game.lcdOutput.framebufferIndex\[2\] vssd1 vssd1 vccd1 vccd1
+ net131 sky130_fd_sc_hd__buf_2
Xfanout120 _3181_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
Xfanout142 _0643_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
Xfanout153 net157 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_2
Xfanout164 _0644_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout175 net178 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
XANTENNA__9271__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6212__A1 _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7714__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6346__A allocation.game.collision.dinoY\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5870_ _1792_ _1793_ _1794_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__nand3_1
X_4821_ _0739_ _0745_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_4752_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7540_ _3032_ _3070_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4683_ net229 net227 vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nor2_1
X_7471_ net246 _3086_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6422_ allocation.game.game.score\[3\] _2323_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__and2_1
X_9210_ _0148_ _0407_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9141_ clknet_leaf_17_clk _0205_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6353_ _2276_ _2237_ _2272_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__and3b_1
X_5304_ _1222_ _1225_ _1226_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21o_1
X_9072_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[18\] net189 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6284_ allocation.game.controller.drawBlock.counter\[1\] _2208_ vssd1 vssd1 vccd1
+ vccd1 _2209_ sky130_fd_sc_hd__xnor2_1
X_8023_ _3531_ _3532_ vssd1 vssd1 vccd1 vccd1 _3533_ sky130_fd_sc_hd__and2_1
X_5235_ _1150_ _1157_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9294__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5166_ _1076_ _1090_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__and2b_1
X_5097_ _1016_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__xnor2_1
X_8925_ _4314_ _4323_ _4315_ vssd1 vssd1 vccd1 vccd1 _4375_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_17_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8856_ net266 net40 vssd1 vssd1 vccd1 vccd1 _4306_ sky130_fd_sc_hd__nor2_1
X_7807_ _3317_ _3366_ vssd1 vssd1 vccd1 vccd1 _3369_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8787_ _4222_ _4236_ net44 vssd1 vssd1 vccd1 vccd1 _4237_ sky130_fd_sc_hd__a21o_1
X_5999_ _1819_ _1862_ _1861_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7738_ net51 _3295_ vssd1 vssd1 vccd1 vccd1 _3300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9075__Q allocation.game.dinoJump.dinoMovement vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9408_ clknet_leaf_17_clk _0318_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_7669_ allocation.game.lcdOutput.framebufferIndex\[7\] _3222_ net50 _3220_ vssd1
+ vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9339_ clknet_leaf_5_clk _0019_ net173 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.slow_clk
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold9 _0241_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_2_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4995__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5245__A _1052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5020_ _0943_ _0944_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8661__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_2_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6971_ _2717_ _2718_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__nor2_1
X_8710_ net98 _4155_ _4158_ net76 vssd1 vssd1 vccd1 vccd1 _4161_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5922_ _1843_ _1844_ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5853_ _0762_ net102 vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__nor2_1
X_8641_ net49 _3595_ vssd1 vssd1 vccd1 vccd1 _4092_ sky130_fd_sc_hd__xnor2_1
X_4804_ _0709_ _0727_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__or2_2
X_5784_ _1706_ _1708_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__xnor2_1
X_8572_ _4006_ _4022_ vssd1 vssd1 vccd1 vccd1 _4023_ sky130_fd_sc_hd__nor2_1
X_4735_ _0657_ _0660_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__nor2_1
X_7523_ net251 net248 _3048_ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout216_A allocation.game.cactus1size.clock_div_inst0.reset vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4666_ _0588_ _0595_ _0587_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__a21o_2
XFILLER_0_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7454_ allocation.game.lcdOutput.r_floor _3069_ _3070_ vssd1 vssd1 vccd1 vccd1 _3071_
+ sky130_fd_sc_hd__or3_1
X_4597_ _0530_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoY\[1\] sky130_fd_sc_hd__inv_2
X_7385_ _3011_ allocation.game.cactusMove.x_dist\[5\] _2973_ vssd1 vssd1 vccd1 vccd1
+ _0213_ sky130_fd_sc_hd__mux2_1
X_6405_ allocation.game.game.score\[6\] allocation.game.game.score\[5\] _2321_ _2319_
+ vssd1 vssd1 vccd1 vccd1 _2328_ sky130_fd_sc_hd__a31oi_4
XANTENNA__5155__A _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9124_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[18\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[18\] sky130_fd_sc_hd__dfrtp_1
X_6336_ allocation.game.cactusHeight2\[0\] allocation.game.cactusHeight2\[1\] vssd1
+ vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__xnor2_1
X_9055_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[1\] net189 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[1\] sky130_fd_sc_hd__dfrtp_1
X_6267_ _2065_ _2099_ _2100_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__nand3_1
XANTENNA__8466__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8006_ net427 _3516_ net206 vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__mux2_1
X_5218_ _1124_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__nand2_1
X_6198_ _1480_ _2122_ _1478_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__a21o_1
X_5149_ _1071_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__and2_1
XANTENNA__7612__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8908_ _4319_ _4356_ _4357_ vssd1 vssd1 vccd1 vccd1 _4358_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8839_ _4285_ _4287_ _4288_ _4282_ vssd1 vssd1 vccd1 vccd1 _4289_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5065__A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8159__A1 allocation.game.controller.state\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9000__A _4423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6343__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7906__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7382__A2 _3009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4520_ allocation.game.dinoJump.dinoDelay\[19\] allocation.game.dinoJump.dinoDelay\[20\]
+ allocation.game.dinoJump.dinoDelay\[18\] vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__or3b_1
X_7170_ net237 allocation.game.controller.state\[0\] vssd1 vssd1 vccd1 vccd1 _0000_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6121_ _2045_ _2043_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6052_ _1934_ _1974_ _1973_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__a21o_1
X_5003_ _0926_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__nand2_1
XANTENNA__8398__A1 allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9332__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6954_ _2707_ net91 _2706_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout166_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5905_ _1781_ _1827_ _1826_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9482__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6885_ allocation.game.cactusDist.clock_div_inst1.counter\[10\] _2661_ allocation.game.cactusDist.clock_div_inst1.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8624_ _4068_ _4074_ _4066_ vssd1 vssd1 vccd1 vccd1 _4075_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5836_ _1757_ _1758_ _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_14_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4989__A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8555_ _3999_ _4001_ _4003_ _3997_ vssd1 vssd1 vccd1 vccd1 _4006_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_17_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5767_ _1689_ _1691_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5698_ _0761_ _0887_ _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__and3_1
X_7506_ net355 net53 _3111_ _3118_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__o22a_1
X_8486_ _3268_ _3282_ vssd1 vssd1 vccd1 vccd1 _3939_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_12_Left_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4718_ net164 vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__inv_2
X_4649_ _0577_ _0578_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7437_ allocation.game.lcdOutput.tft.initSeqCounter\[0\] _0430_ vssd1 vssd1 vccd1
+ vccd1 _3054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7368_ _2994_ _3004_ net54 vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7299_ allocation.game.controller.init_module.delay_counter\[14\] allocation.game.controller.init_module.delay_counter\[13\]
+ _2951_ _2954_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__a31o_1
X_9107_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[1\] net183 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__8196__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6319_ _2240_ _2242_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9038_ clknet_leaf_7_clk _0163_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5613__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout79_A _0796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8643__B _3248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4899__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9355__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8553__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7169__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6670_ net225 _2521_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_pixel\[5\]
+ sky130_fd_sc_hd__xor2_1
X_5621_ _1065_ _1534_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8340_ _2295_ net100 _2411_ _3541_ _3633_ vssd1 vssd1 vccd1 vccd1 _3804_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5552_ net61 _1419_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__xnor2_1
X_4503_ allocation.game.controller.drawBlock.idx\[0\] vssd1 vssd1 vccd1 vccd1 _0443_
+ sky130_fd_sc_hd__inv_2
X_8271_ _4456_ net138 vssd1 vssd1 vccd1 vccd1 _3740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5483_ _1390_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__and2_1
X_7222_ allocation.game.dinoJump.count\[13\] allocation.game.dinoJump.count\[12\]
+ allocation.game.dinoJump.count\[14\] _2893_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__and4_1
X_7153_ _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7084_ allocation.game.controller.init_module.idx\[1\] _2758_ _2800_ _2756_ vssd1
+ vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__a31o_1
X_6104_ _2018_ _2028_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6035_ _1959_ _1958_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7986_ net277 net138 vssd1 vssd1 vccd1 vccd1 _3498_ sky130_fd_sc_hd__or2_1
XANTENNA__8791__B2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6937_ allocation.game.scoreCounter.clock_div.counter\[0\] allocation.game.scoreCounter.clock_div.counter\[1\]
+ net91 vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6868_ allocation.game.cactusDist.clock_div_inst1.counter\[4\] _2651_ _2653_ vssd1
+ vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9228__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8607_ _4018_ _4053_ vssd1 vssd1 vccd1 vccd1 _4058_ sky130_fd_sc_hd__nand2_1
X_5819_ _1741_ _1742_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8538_ _3281_ _3947_ _3951_ vssd1 vssd1 vccd1 vccd1 _3990_ sky130_fd_sc_hd__or3_1
XANTENNA__4512__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6799_ _2606_ _2607_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7649__A3 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8469_ net117 _3913_ _3918_ _3921_ vssd1 vssd1 vccd1 vccd1 _3922_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9378__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7034__S net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8654__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9058__RESET_B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7733__A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8829__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6312__A3 _2234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6068__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8564__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7840_ _2973_ _3394_ vssd1 vssd1 vccd1 vccd1 _3395_ sky130_fd_sc_hd__nor2_1
XANTENNA__4673__A_N allocation.game.controller.drawBlock.y_end\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4983_ _0700_ _0701_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__xnor2_4
X_7771_ _3331_ _3332_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__or2_1
XANTENNA__6784__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9510_ net295 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6722_ _2554_ _2555_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9441_ clknet_leaf_15_clk _0350_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6653_ allocation.game.cactusMove.count\[29\] allocation.game.cactusMove.count\[28\]
+ _2507_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9410__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5604_ _1527_ _1528_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__and2_1
X_6584_ _2466_ _2467_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[3\]
+ sky130_fd_sc_hd__nor2_1
X_9372_ clknet_leaf_14_clk _0003_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout129_A allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_8323_ net134 _3523_ _3786_ _3787_ vssd1 vssd1 vccd1 vccd1 _3788_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5535_ net64 _1400_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8254_ _2993_ _3728_ net54 vssd1 vssd1 vccd1 vccd1 _3729_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5466_ _1197_ _1346_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__xor2_1
X_7205_ net84 _2887_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__and2_1
X_8185_ net113 _3673_ _3676_ net100 net205 vssd1 vssd1 vccd1 vccd1 _3677_ sky130_fd_sc_hd__o221a_1
X_5397_ _1272_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7136_ allocation.game.lcdOutput.framebufferIndex\[11\] allocation.game.lcdOutput.framebufferIndex\[10\]
+ _2836_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__and3_1
XANTENNA_input3_A gpio_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7067_ allocation.game.controller.drawBlock.idx\[4\] _2762_ _2763_ vssd1 vssd1 vccd1
+ vccd1 _2787_ sky130_fd_sc_hd__nor3_2
X_6018_ _1941_ _1942_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nand2b_1
X_7969_ _0496_ _0524_ vssd1 vssd1 vccd1 vccd1 _3482_ sky130_fd_sc_hd__xor2_2
XANTENNA__9050__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4546__A_N allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7255__A1 _4459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5520__B _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5320_ _1244_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5251_ _0838_ _1133_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5182_ _1094_ _1102_ _1104_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__nor3_1
XFILLER_0_43_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5711__A _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8941_ net129 _2280_ _4389_ vssd1 vssd1 vccd1 vccd1 _4390_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9073__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8872_ _0401_ net280 _4296_ _4295_ vssd1 vssd1 vccd1 vccd1 _4322_ sky130_fd_sc_hd__a31o_1
X_7823_ _2368_ _3380_ _3381_ vssd1 vssd1 vccd1 vccd1 _3382_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7754_ _2827_ _3283_ _3311_ _3312_ _3315_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__o41a_1
XANTENNA__7638__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4966_ _0705_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_35_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6705_ net441 _2543_ net152 vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4897_ _0819_ _0820_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__xor2_2
X_7685_ _3246_ vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9424_ clknet_leaf_12_clk _0333_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_start\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6636_ allocation.game.cactusMove.count\[21\] allocation.game.cactusMove.count\[22\]
+ _2496_ allocation.game.cactusMove.count\[23\] vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__a31o_1
X_9355_ clknet_leaf_12_clk _0000_ net204 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_6567_ allocation.game.cactusMove.count\[9\] allocation.game.cactusMove.count\[10\]
+ allocation.game.cactusMove.count\[11\] allocation.game.cactusMove.count\[8\] vssd1
+ vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8306_ net273 net137 _3761_ net107 vssd1 vssd1 vccd1 vccd1 _3772_ sky130_fd_sc_hd__a31o_1
X_5518_ net71 _0889_ _1442_ _0918_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__a31o_1
X_6498_ net237 allocation.game.dinoJump.dinoMovement net396 _2408_ vssd1 vssd1 vccd1
+ vccd1 _0010_ sky130_fd_sc_hd__a31o_1
X_9286_ clknet_leaf_1_clk _0101_ net165 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8682__B1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8237_ _3024_ _3029_ vssd1 vssd1 vccd1 vccd1 _3718_ sky130_fd_sc_hd__or2_1
X_5449_ _1372_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__and2_1
X_8168_ net113 net101 _2516_ vssd1 vssd1 vccd1 vccd1 _3662_ sky130_fd_sc_hd__mux2_1
Xfanout110 _0722_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_4
Xfanout121 _0642_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_2
XANTENNA__9416__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 net144 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7119_ net126 _0453_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__or2_1
Xfanout132 allocation.game.lcdOutput.framebufferIndex\[1\] vssd1 vssd1 vccd1 vccd1
+ net132 sky130_fd_sc_hd__clkbuf_2
Xfanout154 net157 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
Xfanout198 net199 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
Xfanout176 net178 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_4
X_8099_ _0654_ _0685_ vssd1 vssd1 vccd1 vccd1 _3602_ sky130_fd_sc_hd__or2_1
X_9513__298 vssd1 vssd1 vccd1 vccd1 _9513__298/HI net298 sky130_fd_sc_hd__conb_1
XANTENNA_fanout61_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8651__B net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4524__X _0462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Left_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9096__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4820_ _0724_ _0743_ _0744_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_32_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _0676_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__nand2_1
X_4682_ allocation.game.cactusMove.cactusMovement net237 vssd1 vssd1 vccd1 vccd1 _0610_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7470_ net249 _3046_ _3073_ _3084_ _3085_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__o311a_1
X_6421_ _2334_ _2342_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9140_ clknet_leaf_18_clk _0204_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.remainingDelayTicks\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4610__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6352_ _0642_ _0662_ _2275_ _2273_ _0661_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__o32a_1
XFILLER_0_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9439__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5303_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__inv_2
X_9071_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[17\] net189 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[17\] sky130_fd_sc_hd__dfrtp_1
X_6283_ _2089_ _2207_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__nor2_1
X_5234_ _1102_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__nor2_1
X_8022_ allocation.game.controller.v\[4\] _3523_ vssd1 vssd1 vccd1 vccd1 _3532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5165_ _1085_ _1088_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout196_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5096_ _1019_ _1020_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__nor2_1
X_8924_ _3275_ _3541_ vssd1 vssd1 vccd1 vccd1 _4374_ sky130_fd_sc_hd__nor2_1
X_8855_ net38 _4304_ _3264_ _4303_ vssd1 vssd1 vccd1 vccd1 _4305_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7806_ net118 _3367_ vssd1 vssd1 vccd1 vccd1 _3368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5998_ _1908_ _1920_ _1921_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout151_X net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8786_ net128 _4212_ _4223_ _4235_ vssd1 vssd1 vccd1 vccd1 _4236_ sky130_fd_sc_hd__a31o_1
XANTENNA__9356__Q allocation.game.controller.state\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4949_ _0823_ _0873_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__or2_1
X_7737_ net50 net48 vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__nand2_1
X_7668_ allocation.game.lcdOutput.framebufferIndex\[6\] _3222_ _3229_ vssd1 vssd1
+ vccd1 vccd1 _3230_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6619_ allocation.game.cactusMove.count\[16\] _2487_ _2489_ _2462_ vssd1 vssd1 vccd1
+ vccd1 allocation.game.cactusMove.n_count\[16\] sky130_fd_sc_hd__o211a_1
X_9407_ clknet_leaf_17_clk _0317_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7599_ allocation.game.cactusDist.lfsr1\[1\] allocation.game.cactusDist.lfsr1\[0\]
+ allocation.game.cactusDist.clock_div_inst0.clk1 vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_42_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9338_ clknet_leaf_6_clk net283 net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9269_ clknet_leaf_2_clk _0061_ net176 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8837__A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6970_ allocation.game.scoreCounter.clock_div.counter\[14\] _2715_ net91 vssd1 vssd1
+ vccd1 vccd1 _2718_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5921_ _0991_ _1845_ _0990_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_0_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_0_clk_X clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9111__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8640_ _4027_ _4050_ _4090_ _4080_ vssd1 vssd1 vccd1 vccd1 _4091_ sky130_fd_sc_hd__or4b_1
X_5852_ _1727_ _1774_ _1775_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__and3_1
X_4803_ _0727_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5783_ _1652_ _1654_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__xnor2_1
X_8571_ net74 _4007_ vssd1 vssd1 vccd1 vccd1 _4022_ sky130_fd_sc_hd__nor2_1
X_4734_ _0648_ _0659_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9497__319 vssd1 vssd1 vccd1 vccd1 net319 _9497__319/LO sky130_fd_sc_hd__conb_1
X_7522_ _3132_ _3020_ _3021_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__or3b_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4665_ _0591_ _0592_ _0590_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__a21o_1
XANTENNA__9261__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7453_ net254 _3019_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__nand2_1
X_4596_ _4457_ net106 _0529_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6404_ _2324_ _2326_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__nand2_1
X_7384_ _3012_ allocation.game.cactusMove.x_dist\[4\] _2973_ vssd1 vssd1 vccd1 vccd1
+ _0212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6335_ _2254_ _2257_ _2258_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__and3b_1
X_9123_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[17\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9054_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[0\] net189 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[0\] sky130_fd_sc_hd__dfrtp_1
X_8005_ net274 net163 _3511_ net241 _3515_ vssd1 vssd1 vccd1 vccd1 _3516_ sky130_fd_sc_hd__a221o_1
X_6266_ allocation.game.controller.drawBlock.counter\[8\] _2189_ vssd1 vssd1 vccd1
+ vccd1 _2191_ sky130_fd_sc_hd__nor2_1
XANTENNA__8466__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5217_ _0843_ _1084_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout199_X net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6197_ _1531_ _2121_ _1529_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__a21o_1
X_5148_ _0791_ _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__and2_1
X_5079_ _1001_ _1003_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__xor2_1
X_8907_ net128 _0466_ _4355_ vssd1 vssd1 vccd1 vccd1 _4357_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8838_ net41 _4283_ vssd1 vssd1 vccd1 vccd1 _4288_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8769_ _4214_ _4218_ vssd1 vssd1 vccd1 vccd1 _4219_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_43_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8340__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9134__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5090__A1 _0731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9284__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7736__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6120_ _2005_ _2033_ _2044_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6051_ _1877_ _1880_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__nand2_1
X_5002_ _0847_ _0850_ _0925_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__nand3_1
X_6953_ allocation.game.scoreCounter.clock_div.counter\[8\] allocation.game.scoreCounter.clock_div.counter\[7\]
+ _2399_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__and3_1
X_5904_ _0778_ _0899_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__nor2_1
X_6884_ allocation.game.cactusDist.clock_div_inst1.counter\[10\] _2661_ _2663_ vssd1
+ vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__o21a_1
X_8623_ net225 net67 _4073_ _4070_ vssd1 vssd1 vccd1 vccd1 _4074_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5835_ _0912_ _1645_ _1759_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout159_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8554_ net220 net99 vssd1 vssd1 vccd1 vccd1 _4005_ sky130_fd_sc_hd__nor2_1
X_5766_ _0901_ _1690_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5697_ net103 _0886_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__nor2_1
X_4717_ net229 allocation.game.cactusMove.x_dist\[2\] vssd1 vssd1 vccd1 vccd1 _0644_
+ sky130_fd_sc_hd__xor2_2
X_8485_ _3891_ _3928_ _3935_ _3937_ vssd1 vssd1 vccd1 vccd1 _3938_ sky130_fd_sc_hd__o211a_1
X_7505_ _0420_ _3115_ _3117_ _3018_ vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__o31a_1
X_4648_ allocation.game.controller.drawBlock.y_end\[6\] allocation.game.controller.drawBlock.y_start\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7436_ _3041_ _3052_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9106_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[0\] net174 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[0\] sky130_fd_sc_hd__dfrtp_1
X_4579_ net264 net106 vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7381__A _3008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7367_ allocation.game.lcdOutput.tft.remainingDelayTicks\[16\] _2993_ net375 vssd1
+ vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__o21ai_1
X_7298_ allocation.game.controller.init_module.delay_counter\[14\] allocation.game.controller.init_module.delay_counter\[13\]
+ net122 vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__o21ai_1
X_6318_ allocation.game.cactusHeight2\[5\] _2239_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__and2_1
X_9037_ clknet_leaf_7_clk _0162_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5613__B _0885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6249_ allocation.game.controller.drawBlock.counter\[17\] _2173_ vssd1 vssd1 vccd1
+ vccd1 _2174_ sky130_fd_sc_hd__nor2_1
XANTENNA__9157__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8077__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 allocation.game.scoreCounter.clock_div.counter\[0\] vssd1 vssd1 vccd1 vccd1
+ net413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__9011__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5620_ _1537_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5551_ net61 _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__nand2_1
X_8270_ _3737_ net145 net233 net153 vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__a2bb2o_1
X_4502_ net126 vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7221_ net448 _2896_ _2898_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5482_ _1387_ _1389_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7152_ _2853_ _2854_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkload13_A clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7083_ allocation.game.controller.init_module.idx\[0\] allocation.game.controller.init_module.idx\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__nand2_1
X_6103_ _2025_ _2026_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6034_ _1916_ _1917_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7985_ net138 _3496_ vssd1 vssd1 vccd1 vccd1 _3497_ sky130_fd_sc_hd__nand2_1
X_6936_ net413 _0019_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8760__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6867_ allocation.game.cactusDist.clock_div_inst1.counter\[4\] _2651_ net159 vssd1
+ vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6798_ net446 _2605_ net153 vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__o21ai_1
X_5818_ _1741_ _1742_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8606_ net47 _4017_ vssd1 vssd1 vccd1 vccd1 _4057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5749_ _1671_ _1672_ _1673_ vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__nand3_1
X_8537_ _3270_ _3988_ vssd1 vssd1 vccd1 vccd1 _3989_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8468_ _3879_ _3914_ _3920_ _3873_ vssd1 vssd1 vccd1 vccd1 _3921_ sky130_fd_sc_hd__o22a_1
X_8399_ _3853_ _3854_ _3842_ vssd1 vssd1 vccd1 vccd1 _3855_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7419_ _3030_ _3037_ allocation.game.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1 vccd1
+ _3038_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_9_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8935__A _0462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8654__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9105__SET_B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9322__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9006__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9472__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4982_ _0700_ _0701_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__xor2_4
X_7770_ _3321_ _3325_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__nor2_1
X_6721_ net453 _2553_ net153 vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9440_ clknet_leaf_10_clk _0349_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.x_start\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_6652_ allocation.game.cactusMove.count\[27\] allocation.game.cactusMove.count\[28\]
+ _2506_ allocation.game.cactusMove.count\[29\] vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9371_ clknet_leaf_13_clk _0002_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5603_ _1052_ _1475_ vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__xnor2_1
X_8322_ _0504_ _3504_ _3512_ _3517_ net134 vssd1 vssd1 vccd1 vccd1 _3787_ sky130_fd_sc_hd__o41a_1
X_6583_ allocation.game.cactusMove.count\[3\] _2465_ net149 vssd1 vssd1 vccd1 vccd1
+ _2467_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_30_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5534_ net65 _1458_ _1456_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__a21oi_1
X_8253_ allocation.game.lcdOutput.tft.remainingDelayTicks\[15\] _2992_ vssd1 vssd1
+ vccd1 vccd1 _3728_ sky130_fd_sc_hd__nand2_1
X_5465_ _1387_ _1389_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__or2_1
X_7204_ allocation.game.dinoJump.count\[9\] _2885_ _2886_ vssd1 vssd1 vccd1 vccd1
+ _2887_ sky130_fd_sc_hd__o21ba_1
X_8184_ _3674_ _3675_ vssd1 vssd1 vccd1 vccd1 _3676_ sky130_fd_sc_hd__nand2_1
X_5396_ _1260_ _1263_ _1271_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nand3_1
XFILLER_0_22_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7135_ allocation.game.lcdOutput.framebufferIndex\[10\] _2836_ vssd1 vssd1 vccd1
+ vccd1 _2838_ sky130_fd_sc_hd__xor2_2
X_7066_ _2770_ _2785_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__nor2_1
X_6017_ _1899_ _1901_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__xnor2_1
X_7968_ net279 net163 net281 vssd1 vssd1 vccd1 vccd1 _3481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7377__Y _3009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7899_ _3430_ _3431_ allocation.game.controller.drawBlock.counter\[9\] net109 vssd1
+ vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__a2bb2o_1
X_6919_ allocation.game.cactusDist.clock_div_inst0.counter\[7\] _2685_ _2687_ vssd1
+ vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9345__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9518__303 vssd1 vssd1 vccd1 vccd1 _9518__303/HI net303 sky130_fd_sc_hd__conb_1
XANTENNA__9495__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5250_ _0831_ _1025_ _1023_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5181_ net60 _1097_ _1099_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__o21bai_1
XANTENNA__8575__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4608__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8940_ net129 _2280_ _2282_ net131 _4388_ vssd1 vssd1 vccd1 vccd1 _4389_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9218__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8871_ _4298_ _4299_ _4313_ _4320_ vssd1 vssd1 vccd1 vccd1 _4321_ sky130_fd_sc_hd__and4bb_1
XANTENNA__8746__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9368__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7822_ _2358_ _2364_ _2367_ _2370_ _2357_ vssd1 vssd1 vccd1 vccd1 _3381_ sky130_fd_sc_hd__a32o_1
X_4965_ _0702_ _0703_ _0704_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7753_ net34 _3314_ vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6704_ allocation.game.cactus1size.clock_div_inst1.counter\[6\] _2543_ vssd1 vssd1
+ vccd1 vccd1 _2544_ sky130_fd_sc_hd__and2_1
XANTENNA__9151__SET_B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout239_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9423_ clknet_leaf_8_clk _0332_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_start\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4896_ _0819_ _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__and2_2
X_7684_ _3222_ _3245_ vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6635_ allocation.game.cactusMove.count\[22\] _2497_ _2499_ vssd1 vssd1 vccd1 vccd1
+ allocation.game.cactusMove.n_count\[22\] sky130_fd_sc_hd__o21a_1
X_9354_ clknet_leaf_11_clk _0286_ net202 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6566_ allocation.game.cactusMove.count\[3\] allocation.game.cactusMove.count\[2\]
+ _2451_ _2452_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__or4_2
X_8305_ _3740_ _3770_ vssd1 vssd1 vccd1 vccd1 _3771_ sky130_fd_sc_hd__nor2_1
X_5517_ net79 _0886_ _0888_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__o21ai_1
X_9285_ clknet_leaf_1_clk _0100_ net166 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6497_ net237 net242 vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8236_ net371 _2988_ vssd1 vssd1 vccd1 vccd1 _3717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5448_ _1319_ _1371_ _1370_ _1366_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__a211o_1
Xfanout122 _2928_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
Xfanout100 _2382_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_4
X_8167_ net414 net206 _3661_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout111 _0640_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
X_5379_ _1300_ _1302_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__xnor2_1
X_8098_ _3597_ _3600_ _3601_ net203 net389 vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__o32a_1
Xfanout133 allocation.game.lcdOutput.framebufferIndex\[1\] vssd1 vssd1 vccd1 vccd1
+ net133 sky130_fd_sc_hd__clkbuf_2
Xfanout144 _0463_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
X_7118_ net126 _0453_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__nand2_1
Xfanout155 net157 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout188 net200 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
X_7049_ allocation.game.controller.drawBlock.idx\[0\] allocation.game.controller.drawBlock.idx\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__or2_1
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
Xfanout177 net178 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_2
Xfanout166 net200 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8673__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8673__B2 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8395__A allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _0649_ net105 vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__or2_1
X_4681_ net237 allocation.game.dinoJump.dinoMovement allocation.game.controller.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_44_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6420_ _2342_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__inv_2
X_6351_ _2274_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__inv_2
X_5302_ _1222_ _1225_ _1226_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__nand3_2
XFILLER_0_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6282_ _0715_ _0895_ net124 net141 vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9070_ clknet_leaf_21_clk allocation.game.dinoJump.next_dinoDelay\[16\] net189 vssd1
+ vssd1 vccd1 vccd1 allocation.game.dinoJump.dinoDelay\[16\] sky130_fd_sc_hd__dfrtp_1
X_5233_ _1096_ _1101_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__and2_1
X_8021_ allocation.game.controller.v\[4\] _3523_ vssd1 vssd1 vccd1 vccd1 _3531_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9040__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5164_ _1085_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__and2b_1
X_5095_ _0857_ _1017_ _1018_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__nor3_1
X_8923_ _4244_ _4372_ vssd1 vssd1 vccd1 vccd1 _4373_ sky130_fd_sc_hd__nand2_1
X_8854_ net258 _0467_ vssd1 vssd1 vccd1 vccd1 _4304_ sky130_fd_sc_hd__xnor2_1
X_7805_ _3300_ _3303_ _3366_ _3365_ net96 vssd1 vssd1 vccd1 vccd1 _3367_ sky130_fd_sc_hd__o32a_1
XFILLER_0_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5997_ _1920_ _1921_ _1908_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__a21oi_1
X_8785_ _4224_ _4234_ vssd1 vssd1 vccd1 vccd1 _4235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4948_ _0871_ _0872_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7736_ net51 _3237_ vssd1 vssd1 vccd1 vccd1 _3298_ sky130_fd_sc_hd__nor2_1
X_4879_ _0793_ net71 vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__nand2_2
X_7667_ allocation.game.lcdOutput.framebufferIndex\[7\] net51 vssd1 vssd1 vccd1 vccd1
+ _3229_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6618_ allocation.game.cactusMove.count\[16\] _2487_ vssd1 vssd1 vccd1 vccd1 _2489_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__4801__A _0710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9406_ clknet_leaf_17_clk _0316_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_7598_ allocation.game.cactusDist.lfsr1\[0\] _3170_ _3171_ vssd1 vssd1 vccd1 vccd1
+ _0268_ sky130_fd_sc_hd__o21ai_1
X_9337_ clknet_leaf_6_clk _0121_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_6549_ allocation.game.dinoJump.dinoDelay\[15\] _2439_ _2415_ vssd1 vssd1 vccd1 vccd1
+ _2442_ sky130_fd_sc_hd__o21ai_1
XANTENNA__8655__A1 _0673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9268_ clknet_leaf_0_clk _0060_ net176 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8219_ allocation.game.lcdOutput.tft.remainingDelayTicks\[3\] _2984_ vssd1 vssd1
+ vccd1 vccd1 _3706_ sky130_fd_sc_hd__nand2_1
X_9199_ _0137_ _0409_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout57_X net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5807__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8894__A1 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9063__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9014__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _0728_ _0741_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7909__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5851_ _1727_ _1775_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__and2_1
X_4802_ _0605_ _0707_ _0708_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5782_ _1706_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__inv_2
X_8570_ net58 _3608_ _4014_ vssd1 vssd1 vccd1 vccd1 _4021_ sky130_fd_sc_hd__or3b_1
X_4733_ _0648_ _0659_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7521_ _0430_ _3061_ _3085_ _3040_ net247 vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9406__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7452_ allocation.game.lcdOutput.r_dino _3066_ allocation.game.lcdOutput.r_cactus
+ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__o21ba_1
X_4664_ _0593_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__inv_2
X_6403_ allocation.game.game.score\[3\] _2323_ allocation.game.game.score\[4\] vssd1
+ vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4595_ _0471_ _0479_ _0528_ net143 vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__a31o_1
X_7383_ allocation.game.cactusMove.x_dist\[2\] _2975_ _3012_ _3013_ vssd1 vssd1 vccd1
+ vccd1 _0211_ sky130_fd_sc_hd__o22a_1
X_6334_ net277 _2256_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__or2_1
X_9122_ clknet_leaf_4_clk allocation.game.cactusMove.n_count\[16\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__8637__A1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9053_ clknet_leaf_9_clk allocation.game.dinoJump.next_dinoY\[7\] net193 vssd1 vssd1
+ vccd1 vccd1 allocation.game.collision.dinoY\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__6648__B1 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7651__B net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6265_ allocation.game.controller.drawBlock.counter\[8\] _2189_ vssd1 vssd1 vccd1
+ vccd1 _2190_ sky130_fd_sc_hd__and2_1
X_8004_ net273 net137 _3505_ _3513_ _3514_ vssd1 vssd1 vccd1 vccd1 _3515_ sky130_fd_sc_hd__o221a_1
X_5216_ _1138_ _1140_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__nand2_1
X_6196_ _2119_ _2120_ _1575_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__a21o_1
X_5147_ _0732_ _0790_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__or2_1
X_5078_ _0938_ _0945_ _0943_ _0841_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8906_ _0466_ _4355_ net128 vssd1 vssd1 vccd1 vccd1 _4356_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8837_ net36 _4281_ vssd1 vssd1 vccd1 vccd1 _4287_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8768_ net268 net267 _4212_ net261 vssd1 vssd1 vccd1 vccd1 _4218_ sky130_fd_sc_hd__a31o_1
XANTENNA__9086__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7719_ net42 net34 _3280_ _3277_ vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_43_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8699_ _3208_ _3672_ vssd1 vssd1 vccd1 vccd1 _4150_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_43_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4531__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9429__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9009__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6050_ _1934_ _1973_ _1974_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__nand3_1
X_5001_ _0847_ _0850_ net60 vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6952_ allocation.game.scoreCounter.clock_div.counter\[7\] allocation.game.scoreCounter.clock_div.counter\[6\]
+ _2398_ allocation.game.scoreCounter.clock_div.counter\[8\] vssd1 vssd1 vccd1 vccd1
+ _2706_ sky130_fd_sc_hd__a31o_1
XANTENNA__9404__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5903_ _1781_ _1826_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__nand3_1
X_6883_ allocation.game.cactusDist.clock_div_inst1.counter\[10\] _2661_ net159 vssd1
+ vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6390__X _2314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8622_ net221 net75 vssd1 vssd1 vccd1 vccd1 _4073_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5834_ _1757_ _1758_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_17_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5765_ _1687_ _1688_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__xnor2_1
X_8553_ net220 net99 vssd1 vssd1 vccd1 vccd1 _4004_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5696_ _0750_ _1620_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__nand2b_1
X_4716_ _0635_ _0636_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__xnor2_1
X_8484_ net39 _3936_ _3929_ _3278_ vssd1 vssd1 vccd1 vccd1 _3937_ sky130_fd_sc_hd__a211o_1
X_7504_ _3056_ _3060_ _3116_ _3114_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__a31o_1
X_4647_ allocation.game.controller.drawBlock.y_start\[6\] allocation.game.controller.drawBlock.y_end\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7435_ net251 allocation.game.lcdOutput.tft.initSeqCounter\[1\] vssd1 vssd1 vccd1
+ vccd1 _3052_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7366_ _2984_ _3003_ net55 vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout107_X net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4578_ _0514_ net106 _0507_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__or3b_1
X_6317_ allocation.game.cactusHeight2\[5\] _2239_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__or2_1
X_9105_ clknet_leaf_3_clk _0201_ net198 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight1\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__7381__B _3009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8477__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7297_ allocation.game.controller.init_module.delay_counter\[13\] _2951_ _2952_ _2953_
+ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9036_ clknet_leaf_7_clk _0161_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_6248_ _1718_ _2116_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_4_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6179_ _2048_ _2103_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_4_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9101__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 allocation.game.controller.init_module.delay_counter\[12\] vssd1 vssd1 vccd1
+ vccd1 net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 allocation.game.controller.drawBlock.x_start\[2\] vssd1 vssd1 vccd1 vccd1
+ net414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9251__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5550_ _1473_ _1474_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4501_ allocation.game.lcdOutput.framebufferIndex\[11\] vssd1 vssd1 vccd1 vccd1 _0441_
+ sky130_fd_sc_hd__inv_2
X_5481_ _1401_ _1404_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__xnor2_1
X_7220_ allocation.game.dinoJump.count\[14\] _2896_ _0472_ vssd1 vssd1 vccd1 vccd1
+ _2898_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8578__A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9470__Q allocation.game.controller.drawBlock.y_end\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6098__A _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7151_ allocation.game.lcdOutput.framebufferIndex\[16\] _2844_ vssd1 vssd1 vccd1
+ vccd1 _2854_ sky130_fd_sc_hd__xor2_1
X_7082_ _2796_ _2799_ _2760_ vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__o21a_1
X_6102_ _2026_ _2025_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6033_ _1954_ _1957_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7984_ _3494_ _3495_ vssd1 vssd1 vccd1 vccd1 _3496_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout171_A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout269_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6935_ net342 _2695_ _2697_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__a21oi_1
X_6866_ _0449_ _2649_ _2652_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6280__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6797_ allocation.game.cactus2size.clock_div_inst1.counter\[9\] _2605_ vssd1 vssd1
+ vccd1 vccd1 _2606_ sky130_fd_sc_hd__and2_1
X_8605_ _4053_ _4055_ _4054_ vssd1 vssd1 vccd1 vccd1 _4056_ sky130_fd_sc_hd__a21oi_1
X_5817_ _0901_ _1690_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_40_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5748_ _0742_ _0887_ _1622_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__a21o_1
X_8536_ _3316_ _3986_ _3987_ _3951_ vssd1 vssd1 vccd1 vccd1 _3988_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5679_ _1578_ _1603_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__and2_1
X_8467_ _3892_ _3919_ _3344_ vssd1 vssd1 vccd1 vccd1 _3920_ sky130_fd_sc_hd__o21ai_1
X_8398_ allocation.game.controller.v\[4\] _3477_ allocation.game.controller.v\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3854_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9124__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7418_ allocation.game.lcdOutput.tft.spi.idle _0428_ net55 vssd1 vssd1 vccd1 vccd1
+ _3037_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7349_ allocation.game.lcdOutput.tft.remainingDelayTicks\[9\] _2988_ vssd1 vssd1
+ vccd1 vccd1 _2989_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9397__RESET_B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9274__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9019_ net254 vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__inv_2
XANTENNA__8935__B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8951__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7838__Y _3393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9006__B _4452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9067__RESET_B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9022__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4981_ _0702_ _0703_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6720_ allocation.game.cactus1size.clock_div_inst1.counter\[12\] _2553_ vssd1 vssd1
+ vccd1 vccd1 _2554_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6651_ allocation.game.cactusMove.count\[28\] _2507_ _2509_ vssd1 vssd1 vccd1 vccd1
+ allocation.game.cactusMove.n_count\[28\] sky130_fd_sc_hd__o21a_1
X_6582_ allocation.game.cactusMove.count\[3\] _2465_ vssd1 vssd1 vccd1 vccd1 _2466_
+ sky130_fd_sc_hd__and2_1
X_9370_ clknet_leaf_13_clk _0001_ net209 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__9147__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5602_ net61 _1525_ _1524_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__a21bo_1
X_8321_ _3504_ _3512_ _3517_ _0504_ vssd1 vssd1 vccd1 vccd1 _3786_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_30_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5533_ _1456_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5725__A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8252_ _3726_ _3727_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__or2_1
X_5464_ _1338_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__nand2_1
X_7203_ allocation.game.dinoJump.count\[9\] net148 _2882_ vssd1 vssd1 vccd1 vccd1
+ _2886_ sky130_fd_sc_hd__and3_1
X_8183_ net224 _2373_ vssd1 vssd1 vccd1 vccd1 _3675_ sky130_fd_sc_hd__nand2_1
X_5395_ _1317_ _1319_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9297__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7134_ _2836_ _2837_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__nor2_1
XANTENNA__8997__B1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7065_ allocation.game.controller.drawBlock.idx\[3\] allocation.game.controller.drawBlock.idx\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__nand2_1
X_6016_ _1937_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout174_X net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7967_ _3475_ net107 net241 vssd1 vssd1 vccd1 vccd1 _3480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6918_ allocation.game.cactusDist.clock_div_inst0.counter\[7\] _2685_ net161 vssd1
+ vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__a21oi_1
X_7898_ allocation.game.controller.drawBlock.counter\[9\] _3427_ net95 vssd1 vssd1
+ vccd1 vccd1 _3431_ sky130_fd_sc_hd__o21ai_1
X_6849_ _2639_ _2640_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__nor2_1
XANTENNA__8921__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9499_ net284 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_8519_ _3967_ _3970_ _3964_ vssd1 vssd1 vccd1 vccd1 _3971_ sky130_fd_sc_hd__a21o_1
XANTENNA__8011__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout87_X net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8681__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8912__B1 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9017__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8856__A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5180_ _1094_ _1102_ _1104_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8870_ _4314_ _4315_ _4318_ vssd1 vssd1 vccd1 vccd1 _4320_ sky130_fd_sc_hd__a21oi_1
X_7821_ _2356_ _3379_ vssd1 vssd1 vccd1 vccd1 _3380_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4768__A1 allocation.game.controller.block_done vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4964_ net79 _0886_ _0888_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__or3_2
X_7752_ _2827_ net42 net40 net37 vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_16_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6703_ net158 _2542_ _2543_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9422_ clknet_leaf_12_clk _0331_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_start\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4895_ _0743_ _0749_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__xnor2_4
X_7683_ allocation.game.lcdOutput.framebufferIndex\[7\] net50 _3240_ vssd1 vssd1 vccd1
+ vccd1 _3245_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout134_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6634_ allocation.game.cactusMove.count\[22\] _2497_ net144 vssd1 vssd1 vccd1 vccd1
+ _2499_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9353_ clknet_leaf_12_clk _0285_ net201 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_6565_ allocation.game.cactusMove.count\[1\] allocation.game.cactusMove.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__or2_1
X_6496_ net238 net77 _2407_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__o21ai_1
X_8304_ net272 _3760_ vssd1 vssd1 vccd1 vccd1 _3770_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9284_ clknet_leaf_1_clk _0099_ net165 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5516_ _0792_ _1440_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8235_ _3034_ _3716_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__or2_1
X_5447_ _1366_ _1370_ _1371_ _1319_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_2_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8766__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout101 _2382_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_2
X_8166_ _0645_ _3502_ _3596_ _3501_ vssd1 vssd1 vccd1 vccd1 _3661_ sky130_fd_sc_hd__a22o_1
Xfanout112 _0640_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5378_ _1251_ _1300_ _1301_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__and3_1
Xfanout123 _2927_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_2
XANTENNA__5190__A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout134 net136 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
X_8097_ _0644_ _0682_ _2406_ _3595_ vssd1 vssd1 vccd1 vccd1 _3601_ sky130_fd_sc_hd__a22o_1
Xfanout145 _0463_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
X_7117_ net130 net126 vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__nand2_1
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dlymetal6s2s_1
X_7048_ allocation.game.controller.init_module.idx\[0\] allocation.game.controller.init_module.idx\[2\]
+ _2758_ _2767_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__o211a_1
Xfanout178 net188 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
Xfanout167 net169 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9312__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout47_A _3248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8999_ _4443_ _4444_ _4447_ vssd1 vssd1 vccd1 vccd1 _4448_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4534__A _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7845__A _3394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8370__A1 _0541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4931__A1 _0797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4709__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7755__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4680_ net282 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus1size.clock_div_inst0.reset
+ sky130_fd_sc_hd__inv_2
XFILLER_0_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6350_ _0635_ _0654_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5301_ net62 _1168_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6281_ net141 _0895_ allocation.game.controller.drawBlock.counter\[0\] vssd1 vssd1
+ vccd1 vccd1 _2206_ sky130_fd_sc_hd__o21ai_1
X_8020_ _0488_ _3528_ _3529_ vssd1 vssd1 vccd1 vccd1 _3530_ sky130_fd_sc_hd__or3_1
X_5232_ _1152_ _1156_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_5_clk clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
X_5163_ _1067_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9335__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5094_ _0857_ _1018_ _1017_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__o21a_1
X_8922_ net261 _3540_ vssd1 vssd1 vccd1 vccd1 _4372_ sky130_fd_sc_hd__or2_1
X_8853_ _0467_ _3811_ vssd1 vssd1 vccd1 vccd1 _4303_ sky130_fd_sc_hd__nor2_1
XANTENNA__9485__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7804_ net99 net74 vssd1 vssd1 vccd1 vccd1 _3366_ sky130_fd_sc_hd__nand2_1
X_5996_ _1874_ _1919_ _1918_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__a21o_1
X_8784_ _4229_ _4233_ _4231_ vssd1 vssd1 vccd1 vccd1 _4234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4947_ net73 _0754_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__or2_1
X_7735_ net56 net50 vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__nand2_2
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4878_ _0710_ _0800_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__nor2_1
X_7666_ _3221_ _3226_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6617_ allocation.game.cactusMove.count\[15\] _2486_ _2488_ _2462_ vssd1 vssd1 vccd1
+ vccd1 allocation.game.cactusMove.n_count\[15\] sky130_fd_sc_hd__o211a_1
XANTENNA__4801__B net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9405_ clknet_leaf_17_clk _0315_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_9336_ clknet_leaf_6_clk _0120_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_7597_ allocation.game.cactusDist.lfsr1\[0\] _3170_ net143 vssd1 vssd1 vccd1 vccd1
+ _3171_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6548_ allocation.game.dinoJump.dinoDelay\[15\] _2439_ vssd1 vssd1 vccd1 vccd1 _2441_
+ sky130_fd_sc_hd__and2_1
X_6479_ allocation.game.scoreCounter.clock_div.counter\[16\] allocation.game.scoreCounter.clock_div.counter\[15\]
+ allocation.game.scoreCounter.clock_div.counter\[14\] _2393_ _2389_ vssd1 vssd1 vccd1
+ vccd1 _2394_ sky130_fd_sc_hd__a41o_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8655__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9267_ clknet_leaf_0_clk _0059_ net179 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_8218_ _0418_ net406 _2515_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9198_ _0136_ _0132_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_8149_ net89 _0676_ vssd1 vssd1 vccd1 vccd1 _3647_ sky130_fd_sc_hd__xor2_2
XANTENNA__7091__B2 allocation.game.controller.drawBlock.y_start\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_29_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9358__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6638__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1__f_clk_X clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7909__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5850_ _1720_ _1726_ _1725_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4801_ _0710_ net80 _0718_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__nor3_2
XFILLER_0_5_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5781_ _1703_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__and2b_1
X_4732_ net121 _0647_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7520_ _3040_ _3085_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9473__Q allocation.game.controller.drawBlock.y_end\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4663_ _0591_ _0592_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__and2_1
X_9503__288 vssd1 vssd1 vccd1 vccd1 _9503__288/HI net288 sky130_fd_sc_hd__conb_1
XFILLER_0_12_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7451_ net254 allocation.game.lcdOutput.r_floor allocation.game.lcdOutput.r_cactus
+ _3018_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__or4_1
X_6402_ allocation.game.game.score\[3\] _2323_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__nor2_1
XANTENNA__7688__A3 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4594_ _0497_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7382_ _3008_ _3009_ _2976_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6333_ net277 _2256_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__nand2_1
X_9121_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[15\] net182 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9052_ clknet_leaf_9_clk allocation.game.dinoJump.next_dinoY\[6\] net193 vssd1 vssd1
+ vccd1 vccd1 allocation.game.collision.dinoY\[6\] sky130_fd_sc_hd__dfstp_1
X_6264_ _2102_ _2104_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__xnor2_1
X_8003_ net107 allocation.game.controller.state\[4\] vssd1 vssd1 vccd1 vccd1 _3514_
+ sky130_fd_sc_hd__and2b_2
X_5215_ _0842_ _1139_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6195_ _1573_ _1574_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__xnor2_1
X_5146_ net73 _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__and2_1
X_5077_ _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__inv_2
XANTENNA__8270__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8905_ net275 _4458_ vssd1 vssd1 vccd1 vccd1 _4355_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8836_ _4285_ vssd1 vssd1 vccd1 vccd1 _4286_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4653__A_N allocation.game.controller.drawBlock.y_start\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5979_ _1902_ _1903_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__nand2_1
XANTENNA__7666__Y _3228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5779__A_N net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8767_ _4214_ _4216_ _4215_ _3970_ _4211_ vssd1 vssd1 vccd1 vccd1 _4217_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_48_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7718_ net126 _3279_ vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_43_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8698_ _4148_ vssd1 vssd1 vccd1 vccd1 _4149_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7649_ allocation.game.lcdOutput.framebufferIndex\[9\] _3204_ net67 _3201_ vssd1
+ vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__a31o_1
X_9319_ clknet_leaf_5_clk _0126_ net174 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9030__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5000_ net64 _0922_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__xor2_1
XANTENNA__8864__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9468__Q allocation.game.controller.drawBlock.y_end\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6951_ net91 _2704_ _2705_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5902_ _0769_ _0903_ _1779_ _1780_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__a22o_1
X_6882_ _2661_ _2662_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__nor2_1
X_8621_ net221 net75 vssd1 vssd1 vccd1 vccd1 _4072_ sky130_fd_sc_hd__xnor2_1
X_5833_ _1702_ _1709_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8552_ net99 _4002_ vssd1 vssd1 vccd1 vccd1 _4003_ sky130_fd_sc_hd__nor2_1
X_5764_ _1688_ _1687_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__nand2b_1
X_7503_ net248 _3112_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__nand2_1
X_5695_ _1584_ _1585_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__xnor2_1
X_4715_ _0634_ _0638_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__xor2_2
X_8483_ _0442_ _0452_ net42 vssd1 vssd1 vccd1 vccd1 _3936_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4646_ allocation.game.controller.drawBlock.y_start\[7\] allocation.game.controller.drawBlock.y_end\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout214_A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7434_ net253 net251 vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4577_ _0486_ _0506_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__nor2_1
X_7365_ net365 _2983_ vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__8758__B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9104_ clknet_leaf_3_clk _0200_ net198 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6316_ allocation.game.cactusHeight2\[5\] _2239_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7296_ allocation.game.controller.init_module.delay_counter\[13\] _2821_ vssd1 vssd1
+ vccd1 vccd1 _2953_ sky130_fd_sc_hd__nor2_1
X_9035_ clknet_leaf_7_clk _0160_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_6247_ _1667_ _2117_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6178_ _2038_ _2047_ _2046_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__a21o_1
XANTENNA__7046__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5129_ _0972_ _1050_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_4_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__9053__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4813__Y _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8819_ _4259_ _4262_ _4268_ vssd1 vssd1 vccd1 vccd1 _4269_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_15_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4542__A _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold92 allocation.game.lcdOutput.tft.spi.counter\[1\] vssd1 vssd1 vccd1 vccd1 net415
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4717__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 allocation.game.cactusDist.clock_div_inst0.counter\[9\] vssd1 vssd1 vccd1
+ vccd1 net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 allocation.game.dinoJump.dinoDelay\[7\] vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__7747__B net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8859__A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4500_ allocation.game.lcdOutput.framebufferIndex\[13\] vssd1 vssd1 vccd1 vccd1 _0440_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_14_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5480_ _1404_ _1401_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__nand2b_1
XANTENNA_1 _0717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8578__B _3256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6098__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7150_ _2845_ _2850_ _2852_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7081_ allocation.game.controller.drawBlock.y_end\[2\] _2779_ _2793_ _2798_ vssd1
+ vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__a211o_1
X_6101_ _1993_ _1994_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__xnor2_1
X_6032_ _1954_ _1955_ _1956_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__nand3_1
XANTENNA__9076__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8776__A1 _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7983_ _0500_ _3492_ vssd1 vssd1 vccd1 vccd1 _3495_ sky130_fd_sc_hd__nand2b_1
XANTENNA__9198__Q allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_6934_ net342 _2695_ net155 vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9509__294 vssd1 vssd1 vccd1 vccd1 _9509__294/HI net294 sky130_fd_sc_hd__conb_1
X_6865_ net159 _2651_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8604_ net227 net52 vssd1 vssd1 vccd1 vccd1 _4055_ sky130_fd_sc_hd__nor2_1
XANTENNA__6280__C _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6796_ net158 _2604_ _2605_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__nor3_1
X_5816_ _1738_ _1740_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5747_ _0762_ net86 vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__nor2_1
X_8535_ _3327_ net70 _3973_ vssd1 vssd1 vccd1 vccd1 _3987_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8466_ net119 net57 vssd1 vssd1 vccd1 vccd1 _3919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7417_ allocation.game.lcdOutput.tft.state\[1\] allocation.game.lcdOutput.tft.state\[0\]
+ _3025_ net401 vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__a31o_1
X_5678_ _1595_ _1601_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__xnor2_1
X_8397_ allocation.game.controller.v\[5\] allocation.game.controller.v\[4\] _3477_
+ vssd1 vssd1 vccd1 vccd1 _3853_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4629_ allocation.game.controller.drawBlock.x_start\[2\] allocation.game.controller.drawBlock.x_end\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__and2b_1
X_7348_ allocation.game.lcdOutput.tft.remainingDelayTicks\[8\] allocation.game.lcdOutput.tft.remainingDelayTicks\[7\]
+ _2987_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_9_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7279_ allocation.game.controller.init_module.delay_counter\[7\] _2941_ vssd1 vssd1
+ vccd1 vccd1 _2942_ sky130_fd_sc_hd__and2_1
XANTENNA__9419__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9018_ net254 vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__inv_2
XANTENNA__8000__A_N net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4789__C1 _0605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8679__A _0673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9099__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6646__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4980_ _0702_ _0703_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__xor2_2
XANTENNA__5278__A _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6650_ allocation.game.cactusMove.count\[28\] _2507_ net145 vssd1 vssd1 vccd1 vccd1
+ _2509_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6581_ _2465_ net147 _2464_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5601_ _1524_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__and2_1
X_8320_ net107 _3781_ _3784_ net241 vssd1 vssd1 vccd1 vccd1 _3785_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_30_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5532_ _1441_ _1454_ _1455_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__nor3_1
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8251_ _3019_ _3032_ _3026_ vssd1 vssd1 vccd1 vccd1 _3727_ sky130_fd_sc_hd__a21oi_1
X_5463_ _0992_ _1337_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__nand2_1
X_7202_ _4460_ _2879_ _2883_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__a21oi_1
X_8182_ net224 _2373_ vssd1 vssd1 vccd1 vccd1 _3674_ sky130_fd_sc_hd__or2_1
X_5394_ _1307_ _1310_ _1317_ _1318_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7249__B2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7249__A1 allocation.game.dinoJump.dinoMovement vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7133_ allocation.game.lcdOutput.framebufferIndex\[9\] _2834_ vssd1 vssd1 vccd1 vccd1
+ _2837_ sky130_fd_sc_hd__nor2_1
XANTENNA__8997__B2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7064_ _2782_ _2783_ allocation.game.controller.drawBlock.idx\[4\] vssd1 vssd1 vccd1
+ vccd1 _2784_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout281_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6015_ _1834_ _1837_ _1937_ _1939_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__a211o_1
X_7966_ _0470_ _3460_ _3477_ vssd1 vssd1 vccd1 vccd1 _3479_ sky130_fd_sc_hd__nor3_2
X_7897_ allocation.game.controller.drawBlock.counter\[9\] _3427_ vssd1 vssd1 vccd1
+ vccd1 _3430_ sky130_fd_sc_hd__and2_1
X_6917_ _2685_ _2686_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6848_ net459 _2638_ net156 vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__o21ai_1
X_8518_ _3969_ vssd1 vssd1 vccd1 vccd1 _3970_ sky130_fd_sc_hd__inv_2
X_6779_ allocation.game.cactus2size.clock_div_inst1.counter\[1\] allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ allocation.game.cactus2size.clock_div_inst1.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2595_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9498_ net320 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8011__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9241__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8449_ _3281_ _3891_ _3901_ _3360_ vssd1 vssd1 vccd1 vccd1 _3902_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__9391__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7820_ _2353_ _2359_ _2384_ _3378_ vssd1 vssd1 vccd1 vccd1 _3379_ sky130_fd_sc_hd__o22a_1
XANTENNA__9114__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4963_ _0707_ _0708_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__xnor2_4
X_7751_ _3312_ vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__inv_2
X_7682_ _3232_ _3243_ vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__or2_1
X_6702_ allocation.game.cactus1size.clock_div_inst1.counter\[5\] allocation.game.cactus1size.clock_div_inst1.counter\[4\]
+ _2539_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9421_ clknet_leaf_12_clk _0330_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_start\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_6633_ _2497_ _2498_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[21\]
+ sky130_fd_sc_hd__nor2_1
X_4894_ _0722_ net72 net80 vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__a21o_2
XANTENNA__9264__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6564_ allocation.game.cactusMove.count\[5\] allocation.game.cactusMove.count\[4\]
+ allocation.game.cactusMove.count\[6\] allocation.game.cactusMove.count\[7\] vssd1
+ vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__or4b_1
XFILLER_0_42_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9352_ clknet_leaf_1_clk _0284_ net165 vssd1 vssd1 vccd1 vccd1 allocation.game.bcd_ones\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout127_A allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6495_ net238 _2381_ net240 vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__o21ai_1
X_8303_ _3767_ _3768_ vssd1 vssd1 vccd1 vccd1 _3769_ sky130_fd_sc_hd__nor2_1
X_9283_ clknet_leaf_1_clk _0098_ net165 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5515_ _1197_ _1393_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__xor2_1
X_8234_ _2988_ _3715_ net54 vssd1 vssd1 vccd1 vccd1 _3716_ sky130_fd_sc_hd__a21oi_1
X_5446_ _1317_ _1318_ _1307_ _1310_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8766__B net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8165_ net480 net206 _3502_ _3660_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__a31o_1
Xfanout113 _0627_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout102 _0906_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5377_ _1251_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__nand2_1
X_7116_ _0695_ _2824_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__nand2_1
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
X_8096_ _3599_ vssd1 vssd1 vccd1 vccd1 _3600_ sky130_fd_sc_hd__inv_2
Xfanout146 net151 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
Xfanout124 _0899_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_4
X_7047_ allocation.game.controller.init_module.idx\[0\] allocation.game.controller.init_module.idx\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__nand2_1
XANTENNA_input1_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout179 net181 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_4
Xfanout157 _2529_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8998_ net104 _3190_ _4104_ _4446_ vssd1 vssd1 vccd1 vccd1 _4447_ sky130_fd_sc_hd__o31a_1
X_7949_ _4456_ _0525_ net138 vssd1 vssd1 vccd1 vccd1 _3463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8022__A allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4931__A2 _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8168__S _2516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9531__313 vssd1 vssd1 vccd1 vccd1 _9531__313/HI net313 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8830__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9137__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9287__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__8361__A2 _0541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4922__A2 _0846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5300_ net62 _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__nand2_1
XANTENNA__6124__A1 _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6280_ allocation.game.controller.drawBlock.counter\[0\] net141 _0895_ vssd1 vssd1
+ vccd1 vccd1 _2205_ sky130_fd_sc_hd__or3_1
X_5231_ _0924_ _1155_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__xnor2_1
X_5162_ _0845_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__nor2_1
X_5093_ _0833_ _0856_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__nor2_1
X_8921_ _4368_ _4370_ net258 _4364_ vssd1 vssd1 vccd1 vccd1 _4371_ sky130_fd_sc_hd__a2bb2o_1
X_8852_ _4294_ _4301_ vssd1 vssd1 vccd1 vccd1 _4302_ sky130_fd_sc_hd__nand2_1
X_8783_ net133 net278 _4232_ vssd1 vssd1 vccd1 vccd1 _4233_ sky130_fd_sc_hd__a21oi_1
X_7803_ _3200_ net68 vssd1 vssd1 vccd1 vccd1 _3365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7946__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5995_ _1874_ _1918_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__nand3_1
X_7734_ _3295_ vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__inv_2
X_4946_ net73 _0754_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4877_ _0709_ net71 vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__nand2_1
X_7665_ _3221_ _3226_ vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6616_ _2487_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__inv_2
X_9404_ clknet_leaf_17_clk _0314_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7596_ net373 allocation.game.cactusDist.lfsr1\[1\] vssd1 vssd1 vccd1 vccd1 _3170_
+ sky130_fd_sc_hd__nand2_1
X_9335_ clknet_leaf_6_clk _0119_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4801__C _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6547_ _2439_ _2440_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6478_ allocation.game.scoreCounter.clock_div.counter\[9\] allocation.game.scoreCounter.clock_div.counter\[8\]
+ allocation.game.scoreCounter.clock_div.counter\[7\] _2391_ vssd1 vssd1 vccd1 vccd1
+ _2393_ sky130_fd_sc_hd__a31o_1
X_9266_ clknet_leaf_2_clk _0058_ net181 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__7863__A1 allocation.game.controller.drawBlock.state\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_8217_ _3699_ _3701_ _3705_ net207 net449 vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__o32a_1
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9197_ _0135_ _0131_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_5429_ _1344_ _1350_ _1352_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__nand3_1
X_8148_ _3638_ _3641_ _3646_ net206 net379 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__o32a_1
XFILLER_0_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4529__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8079_ _3569_ _3574_ _3585_ vssd1 vssd1 vccd1 vccd1 _3586_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4816__Y _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7856__A allocation.game.controller.drawBlock.state\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8304__X _3770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8974__X _4423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6654__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4800_ net80 _0722_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5780_ _1597_ _1704_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__nor2_1
X_4731_ net121 _0647_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4662_ allocation.game.controller.drawBlock.y_start\[1\] allocation.game.controller.drawBlock.y_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7450_ allocation.game.lcdOutput.r_dino _3066_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6401_ allocation.game.game.score\[3\] allocation.game.game.score\[4\] _2323_ vssd1
+ vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4593_ net280 allocation.game.controller.v\[0\] _0496_ vssd1 vssd1 vccd1 vccd1 _0527_
+ sky130_fd_sc_hd__a21oi_1
X_9120_ clknet_leaf_5_clk allocation.game.cactusMove.n_count\[14\] net184 vssd1 vssd1
+ vccd1 vccd1 allocation.game.cactusMove.count\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7381_ _3008_ _3009_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6332_ _0437_ _2255_ _2238_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__o21a_1
XANTENNA__9302__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9051_ clknet_leaf_3_clk allocation.game.dinoJump.next_dinoY\[5\] net193 vssd1 vssd1
+ vccd1 vccd1 allocation.game.collision.dinoY\[5\] sky130_fd_sc_hd__dfstp_1
X_6263_ _2042_ _2105_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8002_ _3494_ _3503_ _3512_ vssd1 vssd1 vccd1 vccd1 _3513_ sky130_fd_sc_hd__a21o_1
X_5214_ _1135_ _1137_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6194_ _1617_ _2118_ _1615_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout194_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5145_ _1067_ _1069_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5076_ _0999_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__or2_1
XANTENNA__5084__B2 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8904_ net275 _3522_ _4352_ vssd1 vssd1 vccd1 vccd1 _4354_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_46_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8835_ net41 _4283_ _4284_ net44 vssd1 vssd1 vccd1 vccd1 _4285_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5978_ _1851_ _1852_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__xnor2_1
X_8766_ net259 net37 vssd1 vssd1 vccd1 vccd1 _4216_ sky130_fd_sc_hd__nor2_2
X_4929_ _0732_ _0790_ _0828_ _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_47_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8697_ _0657_ _3228_ vssd1 vssd1 vccd1 vccd1 _4148_ sky130_fd_sc_hd__xnor2_1
X_7717_ net132 net130 vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8325__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7648_ allocation.game.lcdOutput.framebufferIndex\[9\] net66 vssd1 vssd1 vccd1 vccd1
+ _3210_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7579_ allocation.game.cactus1size.clock_div_inst1.clk1 allocation.game.cactus1size.lfsr2\[0\]
+ allocation.game.cactus1size.lfsr2\[1\] net143 vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__a31o_1
X_9318_ clknet_leaf_5_clk _0125_ net172 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8300__A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9249_ clknet_leaf_0_clk _0070_ net176 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8494__D1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout62_X net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9325__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__9475__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6950_ allocation.game.scoreCounter.clock_div.counter\[7\] _2399_ vssd1 vssd1 vccd1
+ vccd1 _2705_ sky130_fd_sc_hd__or2_1
X_5901_ _1823_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6881_ net485 _2660_ net152 vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8620_ _4069_ _4070_ _4061_ _4062_ vssd1 vssd1 vccd1 vccd1 _4071_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _1751_ _1754_ _1755_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_17_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5763_ _0914_ _1637_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__xnor2_1
X_8551_ net221 net220 _3674_ vssd1 vssd1 vccd1 vccd1 _4002_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4714_ net111 vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7502_ net250 _3041_ _3074_ _3079_ _3094_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__o2111a_1
X_5694_ net72 _0746_ _1618_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__and3_1
X_8482_ _3917_ _3934_ vssd1 vssd1 vccd1 vccd1 _3935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4645_ _0572_ _0573_ _0543_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7433_ net253 net251 vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout207_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4576_ _0513_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoY\[6\] sky130_fd_sc_hd__inv_2
X_7364_ _2983_ _3002_ net55 vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8758__C net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9103_ clknet_leaf_3_clk _0199_ net195 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight1\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_6315_ allocation.game.cactusHeight2\[3\] allocation.game.cactusHeight2\[4\] _2238_
+ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7295_ net403 _2949_ _2952_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__o21a_1
X_9034_ clknet_leaf_7_clk _0159_ net187 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6246_ allocation.game.controller.drawBlock.counter\[19\] _2170_ vssd1 vssd1 vccd1
+ vccd1 _2171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6575__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6177_ _2052_ _2053_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_4_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5128_ _0897_ _0915_ _0912_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_49_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ _0982_ _0975_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_28_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4823__A _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8818_ net41 _4256_ vssd1 vssd1 vccd1 vccd1 _4268_ sky130_fd_sc_hd__nand2_1
XANTENNA__9348__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8749_ _4092_ _4093_ vssd1 vssd1 vccd1 vccd1 _4200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8030__A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7809__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold82 allocation.game.controller.drawBlock.y_start\[5\] vssd1 vssd1 vccd1 vccd1
+ net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 allocation.game.controller.drawBlock.x_start\[7\] vssd1 vssd1 vccd1 vccd1
+ net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 allocation.game.cactus2size.clock_div_inst1.counter\[1\] vssd1 vssd1 vccd1
+ vccd1 net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 allocation.game.dinoJump.count\[4\] vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8170__A0 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6100_ _2023_ _2024_ _2022_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7080_ net236 _2797_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6031_ _1912_ _1953_ _1952_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__9479__Q allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7982_ _3492_ _3493_ vssd1 vssd1 vccd1 vccd1 _3494_ sky130_fd_sc_hd__or2_1
X_6933_ _2695_ _2696_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8741__A1_N net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5739__A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6864_ _0449_ _2649_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5815_ _0901_ _1738_ _1739_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8603_ net226 net59 vssd1 vssd1 vccd1 vccd1 _4054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6795_ allocation.game.cactus2size.clock_div_inst1.counter\[7\] allocation.game.cactus2size.clock_div_inst1.counter\[8\]
+ _2601_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_40_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5746_ net103 _0888_ _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__or3_1
X_8534_ _3310_ _3904_ _3971_ vssd1 vssd1 vccd1 vccd1 _3986_ sky130_fd_sc_hd__a21oi_1
X_8465_ _3288_ _3322_ _3868_ _3917_ vssd1 vssd1 vccd1 vccd1 _3918_ sky130_fd_sc_hd__a31oi_1
X_5677_ _1595_ _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__and2b_1
X_4628_ _0556_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_26_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7416_ _3020_ _3026_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__or2_1
X_8396_ _3842_ _3852_ _3851_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4559_ net280 allocation.game.controller.v\[0\] _0496_ vssd1 vssd1 vccd1 vccd1 _0497_
+ sky130_fd_sc_hd__and3_1
X_7347_ allocation.game.lcdOutput.tft.remainingDelayTicks\[6\] _2986_ vssd1 vssd1
+ vccd1 vccd1 _2987_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7278_ net123 _2940_ _2941_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_38_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6229_ _2137_ _2153_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__xnor2_1
X_9017_ net254 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__inv_2
XANTENNA__8216__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5649__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5450__A1 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5559__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6580_ allocation.game.cactusMove.count\[1\] allocation.game.cactusMove.count\[0\]
+ allocation.game.cactusMove.count\[2\] vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5600_ _1471_ _1523_ _1522_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5531_ _1441_ _1454_ _1455_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8250_ _2992_ _3725_ net54 vssd1 vssd1 vccd1 vccd1 _3726_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7201_ net150 _2884_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5462_ _0731_ _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__nand2_1
XANTENNA__9043__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8181_ _0622_ _2311_ vssd1 vssd1 vccd1 vccd1 _3673_ sky130_fd_sc_hd__nor2_1
X_5393_ _1266_ _1316_ _1315_ _1296_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7132_ allocation.game.lcdOutput.framebufferIndex\[9\] _2834_ vssd1 vssd1 vccd1 vccd1
+ _2836_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7063_ allocation.game.controller.drawBlock.idx\[1\] _2771_ allocation.game.controller.drawBlock.x_end\[8\]
+ allocation.game.controller.drawBlock.idx\[0\] vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__and4bb_1
XANTENNA__4909__Y _0834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload11_A clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6014_ _1895_ _1936_ _1935_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7965_ _3477_ vssd1 vssd1 vccd1 vccd1 _3478_ sky130_fd_sc_hd__inv_2
X_7896_ net94 _3428_ _3429_ net108 allocation.game.controller.drawBlock.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__a32o_1
X_6916_ net456 _2683_ net155 vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6847_ allocation.game.cactus2size.clock_div_inst0.counter\[12\] _2638_ vssd1 vssd1
+ vccd1 vccd1 _2639_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6778_ allocation.game.cactus2size.clock_div_inst1.counter\[1\] allocation.game.cactus2size.clock_div_inst1.counter\[0\]
+ allocation.game.cactus2size.clock_div_inst1.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2594_ sky130_fd_sc_hd__nand3_1
XFILLER_0_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5729_ _1599_ _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__and2_1
X_8517_ net56 _3298_ net70 _3968_ vssd1 vssd1 vccd1 vccd1 _3969_ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9497_ net319 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XANTENNA__8685__A1 _3208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8448_ net114 _3899_ _3900_ _3894_ vssd1 vssd1 vccd1 vccd1 _3901_ sky130_fd_sc_hd__a31o_1
X_8379_ _0512_ allocation.game.dinoJump.next_dinoY\[7\] _3839_ vssd1 vssd1 vccd1 vccd1
+ _3840_ sky130_fd_sc_hd__or3b_2
XANTENNA__9066__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__8600__A1 net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4464__Y _0401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ _0707_ _0708_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__xor2_4
X_7750_ allocation.game.lcdOutput.framebufferIndex\[0\] net133 vssd1 vssd1 vccd1 vccd1
+ _3312_ sky130_fd_sc_hd__or2_2
X_4893_ _0792_ _0817_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__xnor2_1
XANTENNA__9409__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7681_ allocation.game.lcdOutput.framebufferIndex\[5\] _3229_ _3239_ vssd1 vssd1
+ vccd1 vccd1 _3243_ sky130_fd_sc_hd__nand3_1
X_6701_ allocation.game.cactus1size.clock_div_inst1.counter\[4\] _2539_ allocation.game.cactus1size.clock_div_inst1.counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9420_ clknet_leaf_8_clk _0329_ vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.y_start\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_6632_ allocation.game.cactusMove.count\[21\] _2496_ net150 vssd1 vssd1 vccd1 vccd1
+ _2498_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9351_ clknet_leaf_4_clk _0283_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.bcd_ones\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6563_ net348 _2448_ _2450_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoDelay\[20\]
+ sky130_fd_sc_hd__a21oi_1
X_8302_ _3493_ _3527_ _3758_ net137 vssd1 vssd1 vccd1 vccd1 _3768_ sky130_fd_sc_hd__a31o_1
X_6494_ net77 vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5514_ _1437_ _1438_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__nor2_1
X_9282_ clknet_leaf_1_clk _0097_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_8233_ allocation.game.lcdOutput.tft.remainingDelayTicks\[7\] _2987_ allocation.game.lcdOutput.tft.remainingDelayTicks\[8\]
+ vssd1 vssd1 vccd1 vccd1 _3715_ sky130_fd_sc_hd__o21ai_1
X_5445_ _1369_ _1367_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__and2b_1
X_8164_ allocation.game.controller.drawBlock.x_start\[1\] net282 vssd1 vssd1 vccd1
+ vccd1 _3660_ sky130_fd_sc_hd__and2_1
X_7115_ allocation.game.controller.init_module.state\[1\] _2826_ vssd1 vssd1 vccd1
+ vccd1 _0399_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout103 _0738_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5376_ _1202_ _1250_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__or2_1
Xfanout136 _3462_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
X_8095_ net113 net101 net230 vssd1 vssd1 vccd1 vccd1 _3599_ sky130_fd_sc_hd__mux2_1
Xfanout147 net151 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
Xfanout125 allocation.game.lcdOutput.framebufferIndex\[14\] vssd1 vssd1 vccd1 vccd1
+ net125 sky130_fd_sc_hd__buf_2
Xfanout114 net116 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_2
X_7046_ net4 allocation.game.lcdOutput.tft.spi.tft_sdi _2760_ _2766_ vssd1 vssd1 vccd1
+ vccd1 net28 sky130_fd_sc_hd__a22o_1
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
Xfanout169 net200 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_2
XANTENNA__6602__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8997_ _4102_ _4107_ _4445_ net116 net89 vssd1 vssd1 vccd1 vccd1 _4446_ sky130_fd_sc_hd__o32a_1
X_7948_ allocation.game.controller.v\[3\] allocation.game.controller.v\[2\] _3460_
+ vssd1 vssd1 vccd1 vccd1 _3462_ sky130_fd_sc_hd__a21o_1
XANTENNA__9089__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7879_ net94 _3416_ _3417_ net108 allocation.game.controller.drawBlock.counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6432__S _2320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5837__A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5230_ _1153_ _1154_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5161_ _0842_ _0844_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__nor2_1
X_5092_ _0809_ _0819_ _0987_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__a21o_1
XANTENNA__7624__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8920_ net36 _4366_ _4367_ net38 _4369_ vssd1 vssd1 vccd1 vccd1 _4370_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9231__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8851_ _4226_ _4300_ _4228_ _4292_ vssd1 vssd1 vccd1 vccd1 _4301_ sky130_fd_sc_hd__or4b_1
X_5994_ _1871_ _1873_ _1872_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__a21o_1
X_8782_ allocation.game.lcdOutput.framebufferIndex\[0\] _4456_ net278 net133 vssd1
+ vssd1 vccd1 vccd1 _4232_ sky130_fd_sc_hd__o22a_1
X_7802_ _3315_ _3343_ _3363_ _3269_ vssd1 vssd1 vccd1 vccd1 _3364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7946__B allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4945_ _0864_ _0869_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__xnor2_1
X_7733_ net46 _3292_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__nand2_2
XFILLER_0_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5747__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4876_ net78 _0799_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__nand2_1
XANTENNA__9381__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8888__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7664_ _3223_ _3225_ vssd1 vssd1 vccd1 vccd1 _3226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6615_ allocation.game.cactusMove.count\[15\] _2486_ vssd1 vssd1 vccd1 vccd1 _2487_
+ sky130_fd_sc_hd__and2_1
X_9403_ clknet_leaf_17_clk _0313_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_7595_ net373 _2674_ _3014_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__mux2_1
X_9334_ clknet_leaf_6_clk _0118_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_6546_ net463 _2437_ net90 vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6477_ allocation.game.scoreCounter.clock_div.counter\[9\] allocation.game.scoreCounter.clock_div.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6578__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7026__X net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9265_ clknet_leaf_0_clk _0057_ net188 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_8216_ net240 _2379_ _3704_ _3703_ _3597_ vssd1 vssd1 vccd1 vccd1 _3705_ sky130_fd_sc_hd__a311o_1
X_9196_ _0134_ _0130_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_5428_ _1344_ _1350_ _1352_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__a21o_1
X_8147_ allocation.game.controller.state\[2\] _0625_ _3642_ _3645_ vssd1 vssd1 vccd1
+ vccd1 _3646_ sky130_fd_sc_hd__a31o_1
X_5359_ _0843_ _0797_ _0978_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__mux2_1
X_8078_ _0541_ _3560_ vssd1 vssd1 vccd1 vccd1 _3585_ sky130_fd_sc_hd__xnor2_1
X_7029_ _0446_ allocation.game.scoreCounter.bcd_tens\[3\] allocation.game.scoreCounter.bcd_tens\[1\]
+ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__a21o_1
XFILLER_0_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4545__B allocation.game.controller.v\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5657__A _0761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8879__A1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9104__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__9254__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8803__B2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4730_ _0646_ _0656_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__and2_2
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4661_ allocation.game.controller.drawBlock.y_end\[0\] allocation.game.controller.drawBlock.y_start\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7380_ _3010_ net257 _2973_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__mux2_1
X_6400_ allocation.game.game.score\[2\] _2320_ _2321_ vssd1 vssd1 vccd1 vccd1 _2323_
+ sky130_fd_sc_hd__or3_1
X_4592_ net233 _0526_ vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.next_dinoY\[0\]
+ sky130_fd_sc_hd__nor2_1
X_6331_ allocation.game.cactusHeight2\[1\] allocation.game.cactusHeight2\[2\] vssd1
+ vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9050_ clknet_leaf_3_clk allocation.game.dinoJump.next_dinoY\[4\] net193 vssd1 vssd1
+ vccd1 vccd1 allocation.game.collision.dinoY\[4\] sky130_fd_sc_hd__dfrtp_1
X_6262_ _2017_ _2106_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8001_ _0490_ _3494_ vssd1 vssd1 vccd1 vccd1 _3512_ sky130_fd_sc_hd__nor2_1
X_5213_ _1137_ _1135_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__nand2b_1
X_6193_ _1667_ _2117_ _1665_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__a21boi_1
X_5144_ _1065_ _1066_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout187_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5075_ _0974_ _0998_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8903_ net264 _4352_ vssd1 vssd1 vccd1 vccd1 _4353_ sky130_fd_sc_hd__xnor2_1
XANTENNA__6281__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8834_ _3522_ _3760_ _4277_ vssd1 vssd1 vccd1 vccd1 _4284_ sky130_fd_sc_hd__o21ai_1
XANTENNA__7676__B net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7781__A1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5977_ _1900_ _1901_ _1898_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__a21o_1
X_8765_ net259 net37 vssd1 vssd1 vccd1 vccd1 _4215_ sky130_fd_sc_hd__nand2_1
X_4928_ _0829_ _0852_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4595__A1 _0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8696_ _3358_ _3362_ _4146_ _3284_ _3272_ vssd1 vssd1 vccd1 vccd1 _4147_ sky130_fd_sc_hd__a2111o_1
X_7716_ net34 _3276_ vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7647_ _3205_ _3207_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4859_ _0740_ _0745_ _0744_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__a21oi_4
XANTENNA__9127__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7578_ allocation.game.cactus1size.clock_div_inst1.clk1 allocation.game.cactus1size.lfsr2\[1\]
+ allocation.game.cactus1size.lfsr2\[0\] vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9317_ clknet_leaf_5_clk _0124_ net173 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6529_ allocation.game.dinoJump.dinoDelay\[7\] allocation.game.dinoJump.dinoDelay\[6\]
+ _2423_ allocation.game.dinoJump.dinoDelay\[8\] vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9248_ clknet_leaf_1_clk _0069_ net176 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8494__C1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9277__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5940__A _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9179_ clknet_leaf_15_clk net332 vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.spi.dataShift\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__8050__X _3559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5900_ net87 _0903_ _1823_ _1824_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__nand4_1
XFILLER_0_15_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6880_ allocation.game.cactusDist.clock_div_inst1.counter\[9\] _2660_ vssd1 vssd1
+ vccd1 vccd1 _2661_ sky130_fd_sc_hd__and2_1
X_5831_ _1754_ _1755_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_17_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7496__B _3066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5762_ _1684_ _1686_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8550_ net221 _3674_ net220 vssd1 vssd1 vccd1 vccd1 _4001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4713_ _0631_ _0639_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__xnor2_1
X_7501_ net248 _3112_ _3113_ _3044_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__o211a_1
X_5693_ _1586_ _1587_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__xor2_1
X_8481_ _3282_ _3341_ _3361_ _3927_ vssd1 vssd1 vccd1 vccd1 _3934_ sky130_fd_sc_hd__a31o_1
XANTENNA__8401__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4644_ _0543_ _0573_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__nand2b_2
X_7432_ _3022_ _3048_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4575_ net233 _0512_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__or2_1
X_7363_ net363 net326 vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__nand2_1
X_7294_ net123 _2951_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__nor2_1
X_9102_ clknet_leaf_9_clk _0198_ net195 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6314_ allocation.game.cactusHeight2\[0\] allocation.game.cactusHeight2\[1\] allocation.game.cactusHeight2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9033_ clknet_leaf_5_clk _0158_ net186 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6245_ _1617_ _2118_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6575__B _2461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6176_ _2065_ _2099_ _2100_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5127_ _0897_ _0915_ _0912_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__o21a_2
X_5058_ _0975_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7687__A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4823__B net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8817_ _4262_ _4266_ vssd1 vssd1 vccd1 vccd1 _4267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8748_ net49 _3595_ vssd1 vssd1 vccd1 vccd1 _4199_ sky130_fd_sc_hd__and2_1
X_8679_ _0673_ _4122_ vssd1 vssd1 vccd1 vccd1 _4130_ sky130_fd_sc_hd__and2_1
XANTENNA__5517__B1 _0888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold50 allocation.game.cactusDist.clock_div_inst0.clk1 vssd1 vssd1 vccd1 vccd1 net373
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 allocation.game.controller.init_module.idx\[3\] vssd1 vssd1 vccd1 vccd1 net384
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 allocation.game.cactusMove.drawDoneCactus vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 _0067_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7868__Y _3410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold94 allocation.game.controller.init_module.delay_counter\[17\] vssd1 vssd1 vccd1
+ vccd1 net417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5845__A _0741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6030_ _0762_ net124 vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__nor2_1
X_7981_ _0495_ _0500_ vssd1 vssd1 vccd1 vccd1 _3493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6932_ net440 _2694_ net155 vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__o21ai_1
X_6863_ net152 _2646_ _2649_ _2650_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5814_ _1686_ _1737_ _1736_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8602_ net226 net59 vssd1 vssd1 vccd1 vccd1 _4053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6794_ allocation.game.cactus2size.clock_div_inst1.counter\[7\] _2601_ allocation.game.cactus2size.clock_div_inst1.counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5745_ _0742_ _0885_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__nand2_1
X_8533_ _3315_ _3960_ _3963_ _3984_ _3343_ vssd1 vssd1 vccd1 vccd1 _3985_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5676_ _1599_ _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__xor2_1
X_8464_ net70 _3870_ _3916_ vssd1 vssd1 vccd1 vccd1 _3917_ sky130_fd_sc_hd__nor3_1
X_4627_ allocation.game.controller.drawBlock.x_end\[3\] allocation.game.controller.drawBlock.x_start\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nand2b_1
X_7415_ allocation.game.lcdOutput.tft.state\[1\] _3026_ _3035_ vssd1 vssd1 vccd1 vccd1
+ _0221_ sky130_fd_sc_hd__a21bo_1
X_8395_ allocation.game.controller.v\[4\] _3477_ vssd1 vssd1 vccd1 vccd1 _3852_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4558_ _0494_ _0495_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7346_ allocation.game.lcdOutput.tft.remainingDelayTicks\[5\] allocation.game.lcdOutput.tft.remainingDelayTicks\[4\]
+ _2985_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__or3_1
X_7277_ allocation.game.controller.init_module.delay_counter\[6\] allocation.game.controller.init_module.delay_counter\[5\]
+ _2937_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_38_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4489_ net247 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__inv_2
X_6228_ _2138_ _2152_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__xnor2_1
X_9016_ net254 vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4818__B _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6159_ _2073_ _2083_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__and2_1
XANTENNA__9315__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__9465__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__8976__A _3181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__8915__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5530_ _1394_ _1395_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5461_ _1382_ _1384_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7200_ allocation.game.dinoJump.count\[8\] _2868_ _2874_ _2878_ vssd1 vssd1 vccd1
+ vccd1 _2884_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8180_ _3670_ _3671_ vssd1 vssd1 vccd1 vccd1 _3672_ sky130_fd_sc_hd__or2_1
X_5392_ _1296_ _1315_ _1316_ _1266_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_23_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7131_ _2834_ _2835_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nor2_1
X_7062_ allocation.game.controller.drawBlock.idx\[3\] _2781_ allocation.game.controller.drawBlock.x_start\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__and3b_1
XANTENNA__9338__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6013_ _1834_ _1837_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7964_ allocation.game.controller.v\[3\] _3476_ vssd1 vssd1 vccd1 vccd1 _3477_ sky130_fd_sc_hd__or2_2
XANTENNA__9488__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
X_6915_ allocation.game.cactusDist.clock_div_inst0.counter\[5\] allocation.game.cactusDist.clock_div_inst0.counter\[6\]
+ _2681_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7895_ allocation.game.controller.drawBlock.counter\[6\] allocation.game.controller.drawBlock.counter\[7\]
+ _3420_ allocation.game.controller.drawBlock.counter\[8\] vssd1 vssd1 vccd1 vccd1
+ _3429_ sky130_fd_sc_hd__a31o_1
X_6846_ net161 _2637_ _2638_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__nor3_1
X_6777_ net394 allocation.game.cactus2size.clock_div_inst1.counter\[0\] _2593_ vssd1
+ vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5728_ _1597_ _1598_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__or2_1
X_8516_ _3237_ _3864_ _3930_ _3873_ vssd1 vssd1 vccd1 vccd1 _3968_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_9496_ net318 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
X_5659_ _0769_ _0892_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__nand2_1
X_8447_ _3895_ _3897_ _3898_ _3371_ vssd1 vssd1 vccd1 vccd1 _3900_ sky130_fd_sc_hd__o22a_1
X_8378_ _0465_ allocation.game.dinoJump.next_dinoY\[5\] allocation.game.dinoJump.next_dinoY\[2\]
+ _3838_ vssd1 vssd1 vccd1 vccd1 _3839_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7329_ allocation.game.cactusMove.drawDoneCactus _2974_ vssd1 vssd1 vccd1 vccd1 _2975_
+ sky130_fd_sc_hd__and2_2
XANTENNA__6448__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4739__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7769__B net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4961_ _0705_ _0706_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__xor2_4
XFILLER_0_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4892_ _0815_ _0816_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__nor2_1
X_7680_ _3233_ _3241_ vssd1 vssd1 vccd1 vccd1 _3242_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6700_ allocation.game.cactus1size.clock_div_inst1.counter\[4\] _2539_ _2541_ vssd1
+ vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6631_ allocation.game.cactusMove.count\[21\] _2496_ vssd1 vssd1 vccd1 vccd1 _2497_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9350_ clknet_leaf_1_clk _0282_ net171 vssd1 vssd1 vccd1 vccd1 allocation.game.bcd_ones\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8301_ _3493_ _3758_ _3527_ vssd1 vssd1 vccd1 vccd1 _3767_ sky130_fd_sc_hd__a21oi_1
X_6562_ net348 _2448_ net90 vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6493_ _0690_ _0693_ allocation.game.controller.state\[7\] vssd1 vssd1 vccd1 vccd1
+ _2405_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5513_ _1426_ _1436_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__and2_1
X_9281_ clknet_leaf_1_clk _0096_ net168 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusDist.clock_div_inst1.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk clknet_1_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
X_8232_ net54 _3714_ _3036_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5444_ _1366_ _1368_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__or2_1
X_8163_ _0694_ _3464_ _3659_ net203 allocation.game.controller.drawBlock.x_start\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__o32a_1
XFILLER_0_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7114_ _0425_ _2800_ _2825_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_35_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout104 _0672_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
X_5375_ _1297_ _1299_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__nand2_1
Xfanout137 _3461_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
X_8094_ _3597_ vssd1 vssd1 vccd1 vccd1 _3598_ sky130_fd_sc_hd__inv_2
Xfanout126 allocation.game.lcdOutput.framebufferIndex\[3\] vssd1 vssd1 vccd1 vccd1
+ net126 sky130_fd_sc_hd__buf_2
XFILLER_0_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout115 net116 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_2
X_7045_ _2764_ _2765_ net236 vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__o21ai_1
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_2
Xfanout159 net162 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8996_ net121 net69 _4101_ vssd1 vssd1 vccd1 vccd1 _4445_ sky130_fd_sc_hd__o21a_1
XANTENNA__7966__Y _3479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7947_ allocation.game.controller.v\[3\] allocation.game.controller.v\[2\] _3460_
+ vssd1 vssd1 vccd1 vccd1 _3461_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7878_ allocation.game.controller.drawBlock.counter\[0\] allocation.game.controller.drawBlock.counter\[1\]
+ allocation.game.controller.drawBlock.counter\[2\] allocation.game.controller.drawBlock.counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _3417_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_34_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6829_ allocation.game.cactus2size.clock_div_inst0.counter\[5\] _2625_ net156 vssd1
+ vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9479_ clknet_leaf_7_clk _0386_ net194 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.v\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6774__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__9033__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5853__A _0762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4469__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _0842_ _1083_ _1082_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5091_ _0797_ _0978_ _0977_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__a21o_2
XANTENNA__9478__RESET_B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8850_ _4231_ _4297_ _4299_ vssd1 vssd1 vccd1 vccd1 _4300_ sky130_fd_sc_hd__or3_1
X_5993_ net87 _0900_ _1917_ _1915_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__a31o_1
X_8781_ _4454_ _4230_ vssd1 vssd1 vccd1 vccd1 _4231_ sky130_fd_sc_hd__xnor2_1
X_7801_ net42 net40 _3282_ _3361_ _3360_ vssd1 vssd1 vccd1 vccd1 _3363_ sky130_fd_sc_hd__a41o_1
XFILLER_0_17_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7946__C allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4944_ _0821_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__xor2_1
XANTENNA__9407__RESET_B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7732_ _3293_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__inv_2
XANTENNA__5747__B net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4875_ net78 _0799_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__and2_2
X_7663_ _3204_ _3224_ vssd1 vssd1 vccd1 vccd1 _3225_ sky130_fd_sc_hd__xor2_1
X_9402_ clknet_leaf_17_clk _0312_ net214 vssd1 vssd1 vccd1 vccd1 allocation.game.controller.drawBlock.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__9060__RESET_B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6614_ _2486_ net149 _2485_ vssd1 vssd1 vccd1 vccd1 allocation.game.cactusMove.n_count\[14\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7594_ allocation.game.cactus1size.clock_div_inst1.clk1 _2535_ _3014_ vssd1 vssd1
+ vccd1 vccd1 _0266_ sky130_fd_sc_hd__mux2_1
X_9333_ clknet_leaf_6_clk _0117_ net170 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6545_ allocation.game.dinoJump.dinoDelay\[13\] allocation.game.dinoJump.dinoDelay\[14\]
+ _2436_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__and3_1
X_9264_ clknet_leaf_0_clk _0056_ net180 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6476_ allocation.game.scoreCounter.clock_div.counter\[12\] allocation.game.scoreCounter.clock_div.counter\[11\]
+ _2390_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8215_ net217 _3692_ vssd1 vssd1 vccd1 vccd1 _3704_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9195_ _0133_ _0401_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.framebufferIndex\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_5427_ _1299_ _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__nand2_1
X_8146_ net239 _3643_ _3644_ net281 vssd1 vssd1 vccd1 vccd1 _3645_ sky130_fd_sc_hd__a31o_1
X_5358_ _0976_ _0989_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__nor2_1
X_8077_ net107 _3583_ net242 vssd1 vssd1 vccd1 vccd1 _3584_ sky130_fd_sc_hd__o21a_1
X_5289_ _1152_ _1156_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__and2_1
X_7028_ allocation.game.scoreCounter.bcd_tens\[0\] _2754_ _0445_ vssd1 vssd1 vccd1
+ vccd1 net22 sky130_fd_sc_hd__o21ai_1
XANTENNA__9056__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8979_ _4425_ _4427_ vssd1 vssd1 vccd1 vccd1 _4428_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_2_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5657__B _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5673__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload8_A clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ allocation.game.controller.drawBlock.y_start\[1\] allocation.game.controller.drawBlock.y_end\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6679__A _2526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4591_ net106 _0525_ _0522_ net235 vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__o211a_1
X_6330_ net272 _2253_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6261_ _0432_ _2185_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__nand2_1
X_8000_ net107 _3508_ _3510_ vssd1 vssd1 vccd1 vccd1 _3511_ sky130_fd_sc_hd__nand3b_1
X_5212_ _1079_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__or2_1
X_6192_ _1718_ _2116_ _1717_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5143_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__inv_2
XANTENNA__9079__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4646__B allocation.game.controller.drawBlock.y_end\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_5074_ _0974_ _0998_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__and2_1
X_8902_ net275 net272 net268 vssd1 vssd1 vccd1 vccd1 _4352_ sky130_fd_sc_hd__o21a_1
XANTENNA__6281__A2 _0895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8833_ net264 _4277_ vssd1 vssd1 vccd1 vccd1 _4283_ sky130_fd_sc_hd__xor2_1
XANTENNA__4662__A allocation.game.controller.drawBlock.y_start\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5976_ _1896_ _1897_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__xnor2_1
X_8764_ _0468_ _4213_ vssd1 vssd1 vccd1 vccd1 _4214_ sky130_fd_sc_hd__or2_1
X_4927_ _0850_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7378__A_N _3009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8695_ net46 _4096_ _4140_ _4145_ vssd1 vssd1 vccd1 vccd1 _4146_ sky130_fd_sc_hd__o31a_1
X_7715_ net34 _3276_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4858_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7646_ _3205_ _3207_ vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_43_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9316_ clknet_leaf_6_clk _0123_ net173 vssd1 vssd1 vccd1 vccd1 allocation.game.scoreCounter.clock_div.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4789_ _0707_ _0708_ _0713_ _0605_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a211oi_1
X_7577_ net143 _3160_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6528_ allocation.game.dinoJump.dinoDelay\[7\] allocation.game.dinoJump.dinoDelay\[8\]
+ _2425_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6459_ net219 _2377_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__and2_1
X_9247_ clknet_leaf_2_clk _0068_ net177 vssd1 vssd1 vccd1 vccd1 allocation.game.cactus2size.clock_div_inst1.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__8494__B1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9178_ clknet_leaf_18_clk _0240_ vssd1 vssd1 vccd1 vccd1 allocation.game.lcdOutput.tft.initSeqCounter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__8003__A_N net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8129_ _0690_ _3628_ allocation.game.controller.state\[7\] vssd1 vssd1 vccd1 vccd1
+ _3629_ sky130_fd_sc_hd__o21a_1
XANTENNA__5940__B _0908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout48_X net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9221__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__9371__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5830_ _1703_ _1705_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_17_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5761_ net71 _0903_ _1684_ _1685_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__nand4_1
XFILLER_0_9_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4712_ _0634_ _0638_ _0632_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__o21a_1
X_8480_ _3929_ _3932_ _3927_ _3928_ vssd1 vssd1 vccd1 vccd1 _3933_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7500_ allocation.game.lcdOutput.tft.initSeqCounter\[3\] _3045_ vssd1 vssd1 vccd1
+ vccd1 _3113_ sky130_fd_sc_hd__nand2_1
X_5692_ _1615_ _1616_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__nand2_1
X_7431_ _3045_ _3046_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__nor2_1
XANTENNA__8712__A1 _3208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4643_ allocation.game.controller.drawBlock.x_start\[8\] _0416_ vssd1 vssd1 vccd1
+ vccd1 _0573_ sky130_fd_sc_hd__nand2_1
X_4574_ net106 _0510_ _0511_ _0482_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7362_ net326 net55 vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__nor2_1
X_7293_ allocation.game.controller.init_module.delay_counter\[12\] _2949_ vssd1 vssd1
+ vccd1 vccd1 _2951_ sky130_fd_sc_hd__and2_1
X_6313_ net112 _0671_ _0673_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__and3_1
X_9101_ clknet_leaf_9_clk _0197_ net195 vssd1 vssd1 vccd1 vccd1 allocation.game.cactusHeight1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9032_ clknet_leaf_5_clk _0157_ net185 vssd1 vssd1 vccd1 vccd1 allocation.game.dinoJump.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6244_ allocation.game.controller.drawBlock.counter\[20\] _2168_ vssd1 vssd1 vccd1
+ vccd1 _2169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6175_ _2052_ _2053_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__xnor2_1
X_5126_ _1050_ _0972_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_4_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5057_ _0980_ _0981_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8816_ _4259_ _4265_ vssd1 vssd1 vccd1 vccd1 _4266_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4568__A2 allocation.game.controller.v\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_8747_ _4179_ _4197_ net57 vssd1 vssd1 vccd1 vccd1 _4198_ sky130_fd_sc_hd__o21a_1
X_5959_ _1820_ _1863_ _1883_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_47_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8678_ _0675_ _4122_ _0669_ vssd1 vssd1 vccd1 vccd1 _4129_ sky130_fd_sc_hd__o21ai_1
XANTENNA__9244__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7629_ _3178_ _3179_ _3183_ _3189_ vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__9394__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 allocation.game.lcdOutput.tft.remainingDelayTicks\[1\] vssd1 vssd1 vccd1 vccd1
+ net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 allocation.game.controller.state\[3\] vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 allocation.game.controller.color\[8\] vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 allocation.game.cactus2size.clock_div_inst0.clk1 vssd1 vssd1 vccd1 vccd1 net374
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 allocation.game.controller.drawBlock.y_start\[6\] vssd1 vssd1 vccd1 vccd1
+ net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 allocation.game.cactusMove.pixel\[4\] vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__8942__A1 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5845__B net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6022__A _0716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_clk_A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7980_ _0495_ _0524_ _0493_ vssd1 vssd1 vccd1 vccd1 _3492_ sky130_fd_sc_hd__a21oi_1
XANTENNA__9117__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6931_ allocation.game.cactusDist.clock_div_inst0.counter\[12\] _2694_ vssd1 vssd1
+ vccd1 vccd1 _2695_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6862_ allocation.game.cactusDist.clock_div_inst1.counter\[1\] allocation.game.cactusDist.clock_div_inst1.counter\[0\]
+ allocation.game.cactusDist.clock_div_inst1.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _2650_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5813_ _1686_ _1736_ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__nand3_1
XFILLER_0_9_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8601_ _3358_ _3362_ _4051_ _3284_ _3272_ vssd1 vssd1 vccd1 vccd1 _4052_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_31_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8532_ _3269_ _3983_ _3980_ _3977_ vssd1 vssd1 vccd1 vccd1 _3984_ sky130_fd_sc_hd__a211o_1
XANTENNA__9267__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6793_ allocation.game.cactus2size.clock_div_inst1.counter\[7\] _2601_ _2603_ vssd1
+ vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5744_ _1624_ _1626_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5675_ net65 _1551_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__xnor2_1
X_8463_ net114 _3914_ vssd1 vssd1 vccd1 vccd1 _3916_ sky130_fd_sc_hd__or2_1
X_8394_ allocation.game.controller.v\[4\] net85 vssd1 vssd1 vccd1 vccd1 _3851_ sky130_fd_sc_hd__nand2_1
X_4626_ allocation.game.controller.drawBlock.x_start\[3\] allocation.game.controller.drawBlock.x_end\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7414_ _3029_ _3032_ _3026_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_7345_ allocation.game.lcdOutput.tft.remainingDelayTicks\[3\] _2984_ vssd1 vssd1
+ vccd1 vccd1 _2985_ sky130_fd_sc_hd__or2_1
X_4557_ _4457_ allocation.game.controller.v\[1\] vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7276_ allocation.game.controller.init_module.delay_counter\[5\] _2937_ allocation.game.controller.init_module.delay_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4488_ net256 vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6227_ _2139_ _2151_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__xnor2_1
X_9015_ net255 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__inv_2
X_6158_ _0742_ _0894_ _2072_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__a21o_1
X_5109_ _0993_ _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__xor2_1
X_6089_ _1975_ _1977_ _1976_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__a21o_1
XANTENNA__4789__A2 _0708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5986__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput6 net6 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__clkbuf_4
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5856__A _0769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6926__B1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5460_ _1333_ _1382_ _1383_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5391_ _1248_ _1265_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7130_ allocation.game.lcdOutput.framebufferIndex\[7\] _2832_ allocation.game.lcdOutput.framebufferIndex\[8\]
+ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7061_ allocation.game.controller.drawBlock.idx\[2\] allocation.game.controller.drawBlock.idx\[0\]
+ allocation.game.controller.drawBlock.idx\[1\] vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__and3_1
X_6012_ _1895_ _1935_ _1936_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__and3_1
.ends

