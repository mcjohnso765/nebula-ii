/*
* This is a template for your top level test bench!
* You are responsible for having a test bench for your top
* level design. Otherwise, your design will not be part
* of the tape-out.
*
* Please also include test benches for your team_03_WB
* and team_03_Wrapper modules, if needed to verify
* interfacing with the Wishbone Bus.
*
* The command to run this test bench is:
* make tbsim-source-team_03-team_03
*/

`timescale 1 ns / 1 ps

module team_03_tb();

    ///////////////////////////////////
    // Write your test bench code here!
    ///////////////////////////////////

endmodule