* NGSPICE file created from team_07_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt team_07_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_119_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05903_ _01585_ net122 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__nand2_2
X_09671_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\] _04725_ net1135
+ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a21oi_1
X_06883_ _01615_ _02550_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__nor2_1
XANTENNA__07534__B2 _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05117__B _00828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05834_ _01505_ _01511_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__xor2_1
X_08622_ net455 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08553_ net139 _04005_ _03963_ vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__o21ai_1
X_05765_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07504_ _00759_ _01610_ net100 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_18_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08484_ _03817_ _03898_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05696_ _01318_ _01393_ _01394_ _01408_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07435_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] _03014_
+ net481 vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07366_ net975 _02965_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09105_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ _04342_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__a21o_1
X_06317_ _01970_ _01971_ _01972_ _01992_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__and4_1
XFILLER_0_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07065__A3 _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09036_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04291_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06248_ net456 net180 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ net274 net154 net146 net276 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__o22a_1
Xhold351 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\] vssd1 vssd1 vccd1
+ vccd1 net1031 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold373 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_up vssd1
+ vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[39\]
+ vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold395 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1064 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06576__A2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ net464 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06411__B net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _04866_ _04867_ net966 net234 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_29_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07856__A1_N _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911__655 vssd1 vssd1 vccd1 vccd1 net655 _10911__655/LO sky130_fd_sc_hd__conb_1
XFILLER_0_99_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07082__X _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868__543 vssd1 vssd1 vccd1 vccd1 _10868__543/HI net543 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_103_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10713_ clknet_leaf_60_wb_clk_i _00544_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10644_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[1\]
+ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10575_ clknet_leaf_9_wb_clk_i _00443_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07461__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06602__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07516__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10009_ clknet_leaf_21_wb_clk_i _00006_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05550_ _01259_ _01261_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05481_ _00965_ _01175_ _01193_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07220_ _02864_ _02866_ _02869_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__o31a_1
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07151_ net166 _02033_ _02775_ _02803_ _02773_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06102_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__nor3_1
XFILLER_0_42_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06255__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05689__S0 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05400__B _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07082_ _01618_ net249 _02735_ _02127_ _02734_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a221o_4
XANTENNA__06255__B2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06033_ net195 net181 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__nand2_2
XANTENNA__05510__A_N net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout105 _01691_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06558__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_4
Xfanout127 _01594_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout138 _01648_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_4
Xfanout149 _04869_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_2
X_07984_ _01700_ _01732_ _03375_ _03526_ _03405_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_52_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09723_ net246 _04761_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a21oi_1
X_06935_ _02501_ _02591_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__nor2_1
XANTENNA__07507__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07507__B2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09654_ _04711_ _04712_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__nor2_2
XANTENNA__04967__A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06866_ net283 net430 _02483_ _02536_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_2_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08605_ _01242_ _01248_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05817_ _01496_ _01510_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__nor2_1
X_09585_ _04667_ _04668_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__nor2_1
XANTENNA__06191__B1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06797_ _00696_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02468_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout165_X net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07062__B _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ _03976_ _03990_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__nor2_1
X_05748_ net1091 _01445_ _01447_ _00787_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\]
+ sky130_fd_sc_hd__a22o_1
X_10980__620 vssd1 vssd1 vccd1 vccd1 _10980__620/HI net620 sky130_fd_sc_hd__conb_1
XFILLER_0_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\] _03936_ _03937_
+ _03938_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] vssd1
+ vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o32a_1
X_05679_ _01347_ _01350_ _01366_ _01391_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10108__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07418_ _03004_ _03005_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08398_ _03709_ _03872_ _03850_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05150__X _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07349_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\] vssd1 vssd1
+ vccd1 vccd1 _02958_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05310__B _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ clknet_leaf_3_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[2\]
+ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09019_ net247 _04279_ _04281_ net404 net892 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10291_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[4\]
+ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07077__X _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 _00111_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08113__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] vssd1 vssd1
+ vccd1 vccd1 net850 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06422__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06549__A2 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07237__B _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08067__A_N net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06485__A1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06485__B2 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10627_ clknet_leaf_39_wb_clk_i _00491_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05220__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10558_ clknet_leaf_11_wb_clk_i _00426_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06603__Y _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ clknet_leaf_16_wb_clk_i _00357_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08023__S _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06051__B net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04981_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
XANTENNA__05890__B _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ _01675_ _02021_ net254 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08259__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06651_ _02321_ _02322_ _02323_ _02178_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a31o_1
X_10964__604 vssd1 vssd1 vccd1 vccd1 _10964__604/HI net604 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05602_ net439 net441 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__nand2_2
X_09370_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04530_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__a31o_1
X_06582_ _02196_ _02245_ _02246_ net84 _02255_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a221o_1
X_08321_ _03715_ _03798_ _03752_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_75_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05533_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\]
+ net418 _01206_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08252_ _01281_ _01303_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__nand2_1
X_05464_ _00966_ _01103_ _01107_ _01112_ _01176_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06507__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07203_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ net446 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08183_ _03655_ _03660_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__or2_2
X_05395_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ _00795_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout125_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07134_ _02785_ _02786_ _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07425__B1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07065_ _01679_ _01904_ _01936_ _02687_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__o41a_1
X_06016_ net178 net170 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_54_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05451__A2 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05784__C _01481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07189__C1 _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06400__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ _03415_ _03521_ _03486_ _03519_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__or4b_1
XFILLER_0_57_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09706_ _04750_ _04751_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\]
+ _04730_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a2bb2o_1
X_06918_ _02512_ _02516_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__nor2_1
X_07898_ _03374_ _03382_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__nor2_1
X_09637_ net962 _04700_ _04701_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a21o_1
X_06849_ net255 _02509_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09568_ net482 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04657_ _04658_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08519_ _03981_ _03982_ vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09499_ _00667_ _04626_ net290 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07664__B1 _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05321__A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06219__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ clknet_leaf_3_wb_clk_i _00303_ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05975__B net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ clknet_leaf_56_wb_clk_i _00283_ net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10274_ clknet_leaf_8_wb_clk_i _00266_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10917__661 vssd1 vssd1 vccd1 vccd1 net661 _10917__661/LO sky130_fd_sc_hd__conb_1
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout491 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_2
XANTENNA__10712__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06046__B _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05180_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00890_ vssd1 vssd1
+ vccd1 vccd1 _00893_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07610__A1_N _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ net442 net772 net242 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07821_ _03371_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__nor2_1
X_07752_ _03303_ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__nand2_1
X_04964_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] vssd1
+ vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06703_ _02066_ _02362_ net83 _02079_ _02236_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a221o_1
XANTENNA__10453__RESET_B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ _01678_ _01903_ _01935_ _03174_ _01905_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a311o_1
X_09422_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] _04567_
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\] vssd1
+ vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a31o_1
XANTENNA__07894__A0 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06634_ _02304_ _02306_ _02178_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09353_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06565_ _02218_ _02225_ _02233_ _02238_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout242_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08304_ _03702_ _03778_ _03779_ _03780_ _03711_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a41o_1
X_05516_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ _01223_ _01228_ _01199_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__a211o_1
X_09284_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06496_ _01620_ net270 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ _03674_ _03712_ _03713_ net474 vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__o211a_1
X_05447_ _01060_ _01089_ _01048_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08166_ _00704_ _03647_ _00703_ vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__o21ai_1
X_05378_ net296 _01083_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07949__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07117_ net96 _02770_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__nand2_1
X_08097_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ _00814_ net475 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07048_ _02363_ _02366_ _02702_ _02697_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__o31a_1
XANTENNA__06621__A1 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _04258_ _04260_ _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10961_ net601 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XANTENNA__06137__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06688__A1 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ net648 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06147__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05986__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06434__X _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__B2 _01615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06612__A1 _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10326_ clknet_leaf_25_wb_clk_i _00044_ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ clknet_leaf_4_wb_clk_i _00249_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10188_ clknet_leaf_75_wb_clk_i net712 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06610__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05226__A _00685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__A1 _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06609__X _02282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06350_ _00710_ net213 net177 _01723_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08971__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05301_ net426 _00999_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06281_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] net130 _01934_ _01938_
+ net256 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05232_ _00899_ _00942_ _00944_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__a21oi_1
X_08020_ net716 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05163_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00876_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08053__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__A3 _01475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05406__A2 _01103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05094_ _00809_ _00818_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__or2_1
X_09971_ clknet_leaf_72_wb_clk_i _00076_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08922_ net234 _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nand2_1
XANTENNA__07159__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ net453 _00706_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ _04187_ vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06520__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07804_ _03351_ _03350_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__nand2b_1
X_08784_ _04139_ _04140_ net192 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__a21oi_1
X_05996_ net133 net122 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__nand2_8
XANTENNA__05136__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ net277 _01105_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04947_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07666_ net126 net141 _02260_ _02768_ _01729_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a32o_1
XANTENNA__07331__A2 _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09405_ net476 _04561_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06617_ _01625_ _02140_ _02289_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07597_ _03152_ _03154_ _03155_ _03151_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__o31a_1
XFILLER_0_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09336_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_138_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06548_ net282 _00748_ _02180_ net85 net261 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a32o_1
XANTENNA__07501__D _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07095__A1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09267_ net363 _04426_ _04464_ net928 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_134_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06479_ _02034_ _02035_ _02038_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a31o_2
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903__568 vssd1 vssd1 vccd1 vccd1 _10903__568/HI net568 sky130_fd_sc_hd__conb_1
X_08218_ net457 _03693_ _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06842__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09198_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ _04369_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08149_ net473 _03634_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08910__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ clknet_leaf_44_wb_clk_i _00149_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08347__A1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09544__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07526__A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10042_ _00062_ _00640_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold30 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\] vssd1
+ vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\] vssd1 vssd1
+ vccd1 vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ team_07_WB.instance_to_wrap.audio vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05333__A1 _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ net550 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__06148__Y _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05884__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07086__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06605__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10309_ clknet_leaf_42_wb_clk_i net797 net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05850_ _01534_ _01537_ _01540_ _01541_ _01536_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__a41o_4
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05781_ _01461_ _01462_ _01463_ _01464_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__and4b_1
X_07520_ _01873_ _02744_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__or2_2
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05243__X _00956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07451_ net451 net409 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__and2_2
XFILLER_0_88_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06521__B1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06402_ _02060_ _02071_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07382_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] _02981_
+ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09121_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ _04355_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06333_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _01631_ _02007_
+ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06264_ net176 _01923_ _01925_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06074__X _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05215_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ _00897_ _00915_ _00927_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__a311o_1
X_08003_ _03552_ _03553_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08026__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold500 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
X_06195_ _01855_ _01872_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__o21ai_1
Xhold511 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout205_A _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05146_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1 vssd1 vccd1 vccd1
+ _00859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09954_ clknet_leaf_82_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[3\]
+ net301 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_38_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05077_ net421 _00694_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[0\] _00675_
+ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ _01405_ net438 net436 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__or3b_1
X_09885_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] _01773_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout195_X net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08836_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] _04142_
+ net926 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07552__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08767_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] net775 net232 vssd1
+ vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__mux2_1
X_05979_ _01647_ _01655_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__o21ai_1
X_07718_ _01590_ _01598_ _01065_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__a21oi_1
X_08698_ _00693_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ _01238_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_64_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07081__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07649_ _03204_ _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ clknet_leaf_18_wb_clk_i _00515_ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_101_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06128__C _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09319_ _00661_ _04500_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10591_ clknet_leaf_36_wb_clk_i _00455_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08116__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05983__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07240__A1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06043__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__07240__B2 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput75 net388 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10025_ clknet_leaf_52_wb_clk_i _00002_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10927_ net576 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_85_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05223__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10858_ net533 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10789_ clknet_leaf_76_wb_clk_i _00610_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05510__Y _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05000_ net12 net11 net14 net13 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__or4_1
XANTENNA__06054__B net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09508__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__A2 _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _02506_ _02508_ net174 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05902_ _01585_ net122 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__and2_1
X_09670_ _01763_ _04712_ _04721_ _04726_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a31o_1
X_06882_ _01608_ _02478_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08621_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net455 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__nand2_1
X_05833_ _01506_ _01520_ _01523_ _01525_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__nand4_2
XFILLER_0_55_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ _03611_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__xor2_1
X_05764_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07503_ _03058_ _03061_ _03062_ _03050_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stageDetect
+ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_18_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08483_ net466 net473 _03640_ _03659_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_18_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05695_ net489 _01404_ _01407_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout155_A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07434_ _03014_ _03015_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[18\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07365_ _02965_ _02972_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_rs_enable
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout322_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ net208 _04344_ _04345_ net400 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__a32o_1
X_06316_ _01983_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__or2_1
XANTENNA__06245__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07296_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__nand2_1
X_09035_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04291_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06247_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] net171 _01923_ vssd1
+ vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold330 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold341 _00394_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ net276 net146 _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold352 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold363 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05129_ _00837_ _00838_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\] vssd1 vssd1
+ vccd1 vccd1 net1043 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold385 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] vssd1 vssd1
+ vccd1 vccd1 net1054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09937_ net464 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XANTENNA__06411__C net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09868_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _04228_ net258 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _04166_ _04167_ net193 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__a21oi_1
X_09799_ net1034 _04808_ _04819_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ clknet_leaf_68_wb_clk_i _00543_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909__574 vssd1 vssd1 vccd1 vccd1 _10909__574/HI net574 sky130_fd_sc_hd__conb_1
XFILLER_0_49_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10643_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[0\]
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10574_ clknet_leaf_9_wb_clk_i _00442_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05472__B1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08370__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06602__B _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07516__A2 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ clknet_leaf_51_wb_clk_i _00005_ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_59_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07348__A1_N net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05480_ _00964_ _01109_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07150_ net146 net125 _01710_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06101_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\] _01783_
+ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__or2_2
X_07081_ net96 net94 net88 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06032_ net196 net185 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nor2_8
XFILLER_0_112_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06352__X _02027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout106 _01651_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout117 _01608_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08952__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout128 _01594_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_6
X_07983_ net263 _03354_ _03363_ net262 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__o22a_1
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_09722_ _04731_ _04760_ _04762_ _04730_ net1059 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a32o_1
XANTENNA__05128__B team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ net427 _01652_ _01700_ _02503_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_52_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07507__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07183__X _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net1029 _04711_ _04713_ _04715_ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06865_ net279 _02474_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08604_ _01243_ _01758_ _04035_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand4_2
X_05816_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _01486_
+ _01490_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09584_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\] _04665_ net1071
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06191__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06796_ _00695_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02467_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06191__B2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05144__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08535_ _03974_ _03990_ _03978_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__a21o_1
XANTENNA__07062__C _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05747_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout158_X net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08466_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
X_05678_ _01345_ _01378_ _01390_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07417_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] _03003_
+ net230 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07691__B2 _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03804_ _03847_
+ _00727_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ net491 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _02956_
+ _02957_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_row
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_104_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05310__C _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07279_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__inv_2
X_10290_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[3\]
+ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold160 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__dlygate4sd3_1
X_10835__510 vssd1 vssd1 vccd1 vccd1 _10835__510/HI net510 sky130_fd_sc_hd__conb_1
Xhold193 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\] vssd1 vssd1
+ vccd1 vccd1 net862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06706__B1 _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05989__A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10110__D team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07540__Y _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07682__A1 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10626_ clknet_leaf_39_wb_clk_i net885 net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05995__Y _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ clknet_leaf_13_wb_clk_i _00425_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05445__B1 _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10488_ clknet_leaf_11_wb_clk_i _00356_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07198__B1 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__A1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05229__A team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04980_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06650_ _02107_ _02295_ _02308_ _02139_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22oi_1
XANTENNA__06173__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08974__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10578__Q team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05601_ _01300_ _01313_ _01280_ _01297_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06581_ _02231_ _02253_ _02254_ _02248_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ net462 _03784_ _03796_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05532_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01231_ _01244_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a211o_1
XANTENNA__07122__B1 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08251_ _03685_ _03727_ _03728_ _01384_ net459 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07673__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05463_ _01100_ _01105_ _01111_ _01048_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_31_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06507__B _02180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07202_ _02827_ _02844_ _02847_ _01719_ _02853_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[2\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08182_ net472 net470 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05394_ _01000_ _01003_ _01019_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__or3_2
XFILLER_0_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07133_ _02754_ _02773_ _02781_ _02733_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06228__A2 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout118_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ net128 _01904_ _01936_ _02684_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06523__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06015_ net178 net170 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07189__B1 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05139__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07966_ net276 net108 net269 _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o31a_1
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09705_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] _04749_ _04731_
+ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06917_ _02579_ _02586_ _02587_ _02578_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a31o_1
X_07897_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\] _04698_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__and3b_1
X_06848_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ _04657_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04548_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_136_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06779_ net183 _02447_ _02449_ _02450_ _02432_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08518_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ _03979_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07801__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] vssd1
+ vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06467__A2 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07664__A1 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08449_ _03632_ _03662_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nand2_1
XANTENNA__07664__B2 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05321__B _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ clknet_leaf_3_wb_clk_i _00302_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10342_ clknet_leaf_56_wb_clk_i _00282_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05978__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06433__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10273_ clknet_leaf_8_wb_clk_i _00265_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout90_X net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10105__D team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\] vssd1
+ vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_2
X_10987__627 vssd1 vssd1 vccd1 vccd1 _10987__627/HI net627 sky130_fd_sc_hd__conb_1
XFILLER_0_115_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08852__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ clknet_leaf_35_wb_clk_i _00473_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07820_ _03372_ _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__nor2_1
X_07751_ _03304_ _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__or2_1
X_04963_ net53 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06702_ net115 net112 _02148_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07682_ _02699_ _03238_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07343__B1 _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ _04571_ _04573_ _04574_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07902__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06633_ _02119_ _02289_ _02305_ _02165_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__o22a_1
XANTENNA__07894__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04520_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a21oi_1
X_06564_ _02160_ net85 _02214_ _02237_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06518__A _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08303_ _03702_ _03778_ _03779_ _03780_ _03711_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a41oi_1
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05515_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\] team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__nor2_1
X_09283_ _04475_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06495_ _02119_ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout235_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08234_ _00711_ team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__or3b_2
XFILLER_0_7_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05446_ _01086_ _01096_ _01078_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08165_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] _03647_
+ vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_95_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout402_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05377_ _00966_ _01050_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07116_ net273 net86 net93 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ _03600_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ _03594_ vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06082__B1 _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload80 clknet_leaf_47_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_113_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07047_ _02065_ net84 _02692_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__and3_1
XANTENNA__06621__A2 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04264_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__nor4_1
XANTENNA__07582__B1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _01692_ _03319_ _03491_ _03492_ net106 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__o32a_1
XFILLER_0_138_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10960_ net600 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_74_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09619_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] _04688_ vssd1
+ vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__or2_1
XANTENNA__07885__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06688__A2 _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net647 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_97_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07637__A1 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07637__B2 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10163__RESET_B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10102__CLK clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05986__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10325_ clknet_leaf_25_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06612__A2 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ clknet_leaf_4_wb_clk_i _00248_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10187_ clknet_leaf_71_wb_clk_i net692 net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07722__A _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06679__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06338__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07628__A1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05300_ _00996_ _01005_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06280_ _01933_ _01947_ _01953_ _01956_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a31o_1
XFILLER_0_126_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05231_ net447 _00840_ net394 _00832_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__a31o_1
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05162_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00875_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08053__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05093_ _00809_ _00818_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__nor2_1
X_09970_ clknet_leaf_72_wb_clk_i _00075_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08921_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ _04228_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__or4_1
XANTENNA__06801__A _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ net449 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07803_ _01102_ net111 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08783_ _01454_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__nor2_1
X_05995_ net132 net128 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout185_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07734_ net273 _01104_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__nor2_1
X_04946_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1 vssd1 vccd1
+ vccd1 _00686_ sky130_fd_sc_hd__inv_2
XANTENNA__06119__A1 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07665_ _01811_ net164 _03081_ _03222_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ _04560_ _04559_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__mux2_1
X_06616_ _02265_ _02288_ _02272_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07596_ _02082_ _03079_ _03100_ _02744_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_66_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__a21o_1
XANTENNA__07619__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06547_ net261 net84 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09266_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ net363 _04459_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__and4_1
XANTENNA__07095__A2 _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ net184 net178 _02151_ _01684_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_62_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08217_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel _01296_
+ _03694_ _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a2bb2o_1
X_05429_ _01020_ _01053_ _01068_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__a21oi_1
X_09197_ net402 _04375_ _04412_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08148_ net473 _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08079_ _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10110_ clknet_leaf_58_wb_clk_i team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect
+ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.boomGen.boomPixel
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout98_A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08347__A2 _03814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _00061_ _00639_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_101_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07526__B net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05327__A _01039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold42 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold75 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\] vssd1
+ vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\] vssd1
+ vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10943_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs vssd1 vssd1
+ vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10874_ net549 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05333__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05997__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06445__X _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06605__B _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__B2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10308_ clknet_leaf_43_wb_clk_i net734 net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_120_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10239_ clknet_leaf_74_wb_clk_i net702 net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06349__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05780_ _01465_ _01478_ net477 _01422_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07849__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07849__B2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07450_ net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06521__B2 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06401_ _02074_ _02060_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_44_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07381_ _02974_ _02981_ _02982_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[5\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_29_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09120_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ _04355_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06332_ net285 _00754_ net87 net100 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09051_ net248 _04303_ _04304_ net407 net1121 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_13_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06263_ _01649_ _01938_ _01939_ _01934_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08002_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05214_ _00918_ _00926_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08026__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold501 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\] vssd1
+ vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06194_ _01716_ net103 _01873_ _01874_ _01683_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__o311a_1
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold512 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06037__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05145_ _00855_ _00856_ _00857_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout100_A _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09953_ clknet_leaf_80_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[2\]
+ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_05076_ net426 _00695_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _00674_
+ _00799_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_38_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08904_ net1074 _04217_ net259 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__o21a_1
X_09884_ net1103 net151 net149 _04877_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08835_ _04176_ _04177_ net193 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__a21oi_1
X_08766_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] net866 net232 vssd1
+ vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
X_05978_ net159 _01669_ _01664_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_68_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ net143 _01667_ _01743_ _03270_ _03272_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.borderGen.synchronized_rectangle_pixel
+ sky130_fd_sc_hd__a41o_1
X_04929_ net431 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
X_08697_ _00693_ _01238_ _01242_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07081__B net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07648_ net135 net127 _01743_ _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_64_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07579_ _03130_ _03133_ _03134_ _03137_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08905__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09318_ _00661_ net322 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08265__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ clknet_leaf_36_wb_clk_i _00454_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09249_ net228 _04451_ _04452_ net406 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08921__A team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09765__A1 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07096__X _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06441__A _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_37_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10024_ clknet_leaf_33_wb_clk_i net990 net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input30_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06751__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ net575 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_86_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05998__Y _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ net532 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_137_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ clknet_leaf_1_wb_clk_i _00609_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06019__B1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08042__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06351__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10852__527 vssd1 vssd1 vccd1 vccd1 _10852__527/HI net527 sky130_fd_sc_hd__conb_1
X_06950_ net427 _01566_ _02620_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a21o_1
XANTENNA__08977__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05901_ _01579_ _01581_ _01584_ _01587_ _01593_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a41o_2
X_06881_ net117 _02478_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08620_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04046_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__and3_1
X_05832_ _01506_ _01520_ _01523_ _01525_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08551_ net145 _03652_ _03996_ _04004_ vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__o211a_1
X_05763_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_11_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07502_ _02352_ _03060_ _03059_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08482_ net466 _03637_ _03641_ _03819_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05694_ _01402_ _01406_ net434 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07433_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\] _03013_
+ _02984_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07364_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02970_
+ _02971_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__or3b_1
XFILLER_0_31_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09103_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__nand2_1
X_06315_ _01974_ _01984_ _01990_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07295_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout315_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09034_ net248 _04290_ _04292_ net404 net1051 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__a32o_1
X_06246_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] net180 vssd1 vssd1
+ vccd1 vccd1 _01923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold320 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\] vssd1 vssd1
+ vccd1 vccd1 net1000 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ net279 net161 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__nor2_1
Xhold342 team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\] vssd1 vssd1 vccd1
+ vccd1 net1011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold353 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\] vssd1
+ vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__dlygate4sd3_1
X_05128_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__nand2_1
Xhold364 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[38\]
+ vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold386 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_select
+ vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold397 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__dlygate4sd3_1
X_05059_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] _00788_ vssd1
+ vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__or2_1
X_09936_ net464 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
X_09867_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _04228_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_107_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06725__A1_N _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] _01448_
+ _04160_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or3_1
XANTENNA__06194__C1 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ _04818_ _04811_ _04817_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__and3b_1
XANTENNA__06733__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07930__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05605__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ net239 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10711_ clknet_leaf_68_wb_clk_i _00542_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06497__B1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10642_ clknet_leaf_35_wb_clk_i net882 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06436__A _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10573_ clknet_leaf_9_wb_clk_i _00441_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07461__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09738__A1 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06171__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06421__B1 _02080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955__595 vssd1 vssd1 vccd1 vccd1 _10955__595/HI net595 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_127_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ clknet_leaf_32_wb_clk_i net992 net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07714__B _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07730__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06488__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10909_ net574 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_50_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06100_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\] _01782_
+ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07080_ _01619_ _02209_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__nor2_2
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06031_ net154 _01720_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10893__649 vssd1 vssd1 vccd1 vccd1 net649 _10893__649/LO sky130_fd_sc_hd__conb_1
XFILLER_0_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05249__X _00962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06081__A _01762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06412__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout107 _01650_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08952__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10361__SET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout129 _03653_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_4
X_07982_ _03319_ _03480_ _03536_ _03535_ _03493_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__o32a_1
X_09721_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__inv_2
XANTENNA__07905__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06933_ _02479_ _02485_ _02553_ _02557_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a311o_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10104__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _01764_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__nor2_1
X_06864_ _02475_ _02494_ _02530_ _02534_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_2_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05815_ _00713_ _01501_ _01504_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__a21o_1
X_08603_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01197_ net241 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__a21oi_1
X_09583_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ _04665_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06795_ _00695_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02466_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08534_ _03967_ _03974_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05746_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\] _00771_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] vssd1 vssd1 vccd1 vccd1
+ _01446_ sky130_fd_sc_hd__and4bb_1
XANTENNA__06479__B1 _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__A _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ net415 _00676_ net459 vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o21a_1
X_05677_ net443 _01297_ _01372_ _01388_ net439 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07416_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] _03003_
+ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08396_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] _03870_ _03843_
+ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_34_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07691__A2 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ net411 _00711_ _00796_ _01175_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__o41a_1
XFILLER_0_6_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07278_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__and3_1
XANTENNA__05454__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06229_ _01888_ _01898_ _01908_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[1\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold150 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold161 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\] vssd1 vssd1
+ vccd1 vccd1 net830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\] vssd1 vssd1
+ vccd1 vccd1 net841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__04998__X _00735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06954__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07815__A _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ net830 net151 net149 _04899_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__a22o_1
XANTENNA__06706__A1 _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05989__B _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09408__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05070__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10625_ clknet_leaf_39_wb_clk_i _00489_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10556_ clknet_leaf_11_wb_clk_i _00424_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10487_ clknet_leaf_26_wb_clk_i _00355_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07198__A1 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09940__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06173__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05600_ _01307_ _01308_ _01310_ _01312_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06580_ net125 _01642_ _01699_ _02230_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05920__A2 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05531_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\] net418
+ _01231_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ _01206_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07122__B2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08275__B _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08250_ _01384_ _03728_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__nand2_1
XANTENNA__05251__Y _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05462_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right _00963_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up vssd1 vssd1
+ vccd1 vccd1 _01175_ sky130_fd_sc_hd__or4b_4
XFILLER_0_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07201_ _02846_ _02849_ _02850_ _02851_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ net473 net471 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__and2_1
X_05393_ _01056_ _01063_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07132_ _01676_ _01678_ net162 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07063_ _01678_ _01903_ _01935_ _02715_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a41o_1
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05436__B2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858__533 vssd1 vssd1 vccd1 vccd1 _10858__533/HI net533 sky130_fd_sc_hd__conb_1
XANTENNA__06523__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06014_ net194 net170 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05139__B _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06400__A3 _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07965_ _00753_ net108 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout382_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] _04749_ vssd1
+ vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__and2_1
X_06916_ _02496_ _02581_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__or2_1
X_07896_ _01692_ _03378_ _03406_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05155__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _04699_ _04700_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout170_X net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ net428 _02508_ net251 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06778_ net422 _00986_ net198 _00983_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__o211a_1
X_09566_ net410 _01417_ _01476_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__or3_2
XANTENNA__06538__X _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08517_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] _03979_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__a21oi_1
X_05729_ net474 _00796_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09497_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] _00667_
+ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08861__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ net765 _03921_ net129 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _03718_ _03853_ _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__nor3_1
XFILLER_0_74_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05321__C _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10410_ clknet_leaf_3_wb_clk_i _00301_ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_78_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ clknet_leaf_50_wb_clk_i _00281_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08949__A_N net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10272_ clknet_leaf_8_wb_clk_i _00264_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout83_X net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] vssd1 vssd1
+ vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_2
Xfanout471 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\] vssd1
+ vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_2
Xfanout482 net483 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_79_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07104__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ clknet_leaf_35_wb_clk_i _00472_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10539_ clknet_leaf_29_wb_clk_i _00407_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09935__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970__610 vssd1 vssd1 vccd1 vccd1 _10970__610/HI net610 sky130_fd_sc_hd__conb_1
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07040__B1 _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06394__A2 _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04962_ net1088 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
X_07750_ _01083_ net146 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nor2_1
XANTENNA__09868__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06701_ _01699_ _02266_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07681_ _03098_ _03099_ _03144_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07343__A1 _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09420_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ _04567_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a21o_1
X_06632_ _02268_ _02272_ _02288_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ net223 _04522_ _04523_ net395 net1116 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__a32o_1
X_10929__578 vssd1 vssd1 vccd1 vccd1 _10929__578/HI net578 sky130_fd_sc_hd__conb_1
X_06563_ _02153_ _02234_ _02235_ _02236_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06518__B _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08302_ net412 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__nor3_1
X_05514_ net420 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _01226_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__o21ba_1
X_09282_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06494_ _02155_ _02167_ _02153_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07646__A2 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ _03698_ _03711_ net484 vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_99_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05445_ _01011_ _01059_ _01083_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout130_A _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08164_ _03645_ _03647_ vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05376_ net188 _01015_ _01088_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__o21a_1
XANTENNA__06534__A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05409__A1 _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07115_ net277 net88 _01635_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a21oi_2
X_08095_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ _00814_ net475 vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload70 clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__06082__A1 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ _02138_ net84 _02699_ _02700_ _02362_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_73_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload81 clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_12
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__04989__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08997_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ net263 _03414_ _03416_ net262 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06137__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _03433_ _03429_ _03426_ _03425_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ _04666_ _04687_ _04689_ _04664_ net1040 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__a32o_1
X_10890_ net646 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_66_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09549_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[43\]
+ net266 net288 net218 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05332__B _01039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10324_ clknet_leaf_25_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[1\]
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10255_ clknet_leaf_4_wb_clk_i _00247_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ clknet_leaf_71_wb_clk_i net689 net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07573__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08770__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 _04584_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_2
XANTENNA__05226__C _00828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload6_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__B net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07876__A2 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06619__A _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07628__A2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05230_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08045__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05161_ _00873_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05092_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__or3_1
X_10820__495 vssd1 vssd1 vccd1 vccd1 _10820__495/HI net495 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_90_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08920_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06801__B _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08851_ net449 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net453 vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07564__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _01102_ net111 vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__nand2_1
X_05994_ _01654_ net168 _01683_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__a21oi_4
X_08782_ _01455_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__or2_2
X_04945_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1 vccd1 vccd1
+ _00685_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07733_ net273 _01055_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07632__B _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _02069_ _02872_ _03198_ _02040_ _03083_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09403_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ _00813_ _00815_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a22o_1
XANTENNA__05878__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06615_ _02274_ _02279_ _02266_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07595_ _01675_ _03042_ _01671_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_66_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06248__B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09334_ _04313_ net223 _04511_ net395 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06546_ net215 net186 _01665_ _02219_ _01664_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_138_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09265_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ net403 net227 _04463_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__a22o_1
X_06477_ _01699_ _01901_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_62_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ net457 _01380_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a21oi_1
X_05428_ _01135_ _01138_ _01139_ _01140_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__or4b_1
X_09196_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ net325 _04407_ net1002 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a41o_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06264__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ _03627_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__and2_2
X_05359_ net191 _01004_ _01010_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_112_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00820_ net410 vssd1 vssd1
+ vccd1 vccd1 _03592_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07029_ _02335_ _02349_ _02683_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10040_ _00060_ _00638_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06719__B1_N _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07823__A _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 _00114_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _00112_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10942_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1
+ vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06439__A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05869__B2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ net548 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_112_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06818__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07491__B1 _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06294__B2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06461__X _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10307_ clknet_leaf_42_wb_clk_i net757 net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10238_ clknet_leaf_74_wb_clk_i net701 net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08743__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06349__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ clknet_leaf_26_wb_clk_i _00179_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07733__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06400_ net186 _01642_ _02073_ net201 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_44_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] _02979_
+ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06331_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\] team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ _01962_ _02006_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireHighlightDetect
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06355__Y team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09050_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ _04301_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06285__A1 _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06262_ net456 net155 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__nand2_1
XANTENNA__05700__B net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05213_ _00924_ _00925_ _00923_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__or3b_1
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08001_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06193_ net210 _01670_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold502 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05144_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06371__X _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09952_ clknet_leaf_56_wb_clk_i _00067_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_05075_ _00670_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] _00801_
+ _00802_ _00800_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08903_ _01401_ _01405_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__nor2_1
X_09883_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] _01773_ vssd1
+ vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout295_A _03026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08834_ net1016 _04142_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08765_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] net1053 net237 vssd1
+ vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05977_ _01657_ net170 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout462_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07716_ _03114_ _03271_ _03269_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__a21o_1
X_04928_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1 vssd1
+ vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XANTENNA__06259__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _04114_ _04116_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__o21a_1
XANTENNA__05163__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07081__C net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07647_ _01645_ net143 _01741_ net250 vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_64_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07578_ net123 _03135_ _03132_ _02096_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a211o_1
XANTENNA__06546__X _02220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09317_ net225 _04498_ _04500_ net398 net1045 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_81_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06529_ _01712_ _02088_ _02201_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06276__A1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09248_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04449_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09214__A1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09179_ net207 _04398_ _04400_ net403 net1115 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__A _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06579__A2 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__07537__B net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06441__B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__09267__A1_N net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07528__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ clknet_leaf_33_wb_clk_i _00102_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07528__B2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input23_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05344__Y _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10925_ net669 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XANTENNA__07700__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ net531 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10787_ clknet_leaf_1_wb_clk_i _00608_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07545__A2_N _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06019__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07216__B1 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08323__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08964__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09943__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05248__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05900_ _01579_ _01581_ _01584_ _01587_ _01593_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06880_ _01615_ _02550_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__nand2_1
XANTENNA__06727__C1 _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05831_ _00714_ _01509_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_85_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08550_ _03611_ _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__nand2_1
X_05762_ _01459_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] _01460_ vssd1 vssd1
+ vccd1 vccd1 _01461_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07501_ net95 _01631_ _02009_ _00755_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__and4bb_1
X_05693_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\] _01398_ _01400_
+ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\] vssd1 vssd1 vccd1 vccd1
+ _01406_ sky130_fd_sc_hd__a22o_1
X_08481_ net798 _03952_ net129 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07432_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\] _03013_
+ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__and4b_1
XFILLER_0_9_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09102_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06314_ _01989_ _01988_ _01987_ _01986_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__and4b_1
X_07294_ net740 _02919_ _02923_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[8\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09033_ _04291_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__inv_2
X_06245_ net275 _01920_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout308_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold310 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06176_ net175 net117 net109 net182 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__o22a_1
Xhold321 _00103_ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] vssd1 vssd1
+ vccd1 vccd1 net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold343 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] vssd1 vssd1
+ vccd1 vccd1 net1012 sky130_fd_sc_hd__dlygate4sd3_1
X_05127_ _00835_ _00836_ _00837_ _00839_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__o2bb2a_1
Xhold354 _00025_ vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold365 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 net1034 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold376 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold387 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] vssd1 vssd1
+ vccd1 vccd1 net1056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\] vssd1
+ vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06430__A1 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05058_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ _00787_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__and3_1
X_09935_ net464 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09866_ net1072 net258 _04865_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_107_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _01448_ _04160_ net1047 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_29_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _04797_ _04810_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__nor2_1
XANTENNA__06733__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] net1173 net239 vssd1
+ vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_2_0_wb_clk_i_X clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08679_ _04058_ _04073_ _04100_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ clknet_leaf_68_wb_clk_i _00541_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06497__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06717__A _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10641_ clknet_leaf_35_wb_clk_i _00505_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06436__B net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07446__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ clknet_leaf_9_wb_clk_i _00440_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10006_ clknet_leaf_32_wb_clk_i _00026_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07921__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10210__Q team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06488__A1 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10908_ net573 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XANTENNA__07685__B1 _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10839_ net514 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_67_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09938__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05250__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06030_ net155 _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_1
XANTENNA__09729__A2 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06362__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06412__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 net109 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_4
X_07981_ _01692_ _03475_ _03473_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08952__A3 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] _04754_ vssd1 vssd1
+ vccd1 vccd1 _04761_ sky130_fd_sc_hd__and4_1
XANTENNA__07464__Y _03033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06932_ _02543_ _02554_ _02549_ _02551_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_52_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09362__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05426__A1_N _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06176__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06863_ net117 _02471_ _02531_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07912__A1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08602_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\] _04034_
+ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__and2_1
X_05814_ _00713_ _01501_ _01504_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a21oi_1
X_09582_ _04666_ _04664_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05923__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06794_ net90 _02409_ _02413_ _02438_ _02465_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect
+ sky130_fd_sc_hd__o311a_1
XANTENNA__07480__X _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ _03977_ _03990_ _03991_ _03989_ vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05745_ _01443_ _01445_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_89_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout160_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05712__Y _01425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07676__B1 _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ net460 _03934_ _03935_ net416 _00731_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o221a_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05676_ net439 _01323_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__nand2_1
X_07415_ _03003_ net230 _03002_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[11\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08395_ _01253_ _03733_ _03869_ net458 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_34_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06256__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07346_ _00965_ _02953_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07277_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ _02909_ _02912_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[14\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06543__Y _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__B net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07368__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09016_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04274_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a21o_1
X_06228_ _01738_ _01743_ _01899_ _01900_ _01907_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06159_ net182 _01804_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_76_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold140 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A3 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold151 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold162 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold173 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] vssd1 vssd1
+ vccd1 vccd1 net842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[38\]
+ vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold195 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _01782_ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07815__B _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04850_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06706__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07831__A _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06447__A _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05989__C net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10624_ clknet_leaf_39_wb_clk_i _00488_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10555_ clknet_leaf_11_wb_clk_i _00423_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06642__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486_ clknet_leaf_26_wb_clk_i _00354_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05245__B _00946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05530_ _01197_ _01241_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__or2_1
XANTENNA__06357__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07122__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05461_ _01047_ _01173_ _00964_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07200_ _02040_ _02758_ _02836_ _02848_ _02761_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05392_ _00669_ net393 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__nand2_2
X_08180_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] _00704_
+ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07131_ net137 net105 net162 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07062_ net121 _01903_ _01935_ _02716_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__and4_1
XANTENNA__06633__A1 _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06013_ _01641_ _01674_ _01696_ _01705_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\]
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_11_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07189__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07964_ net133 _03307_ _03487_ _03490_ _03293_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__o311a_1
XFILLER_0_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ net246 _04749_ _04748_ _04733_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a211oi_1
X_06915_ net106 _02497_ _02581_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__or3_1
XANTENNA__06149__B1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ _03448_ _03449_ _03335_ _03440_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__or4bb_1
X_09634_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] _04698_ vssd1
+ vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nand2_1
XANTENNA__05155__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ _02513_ _02516_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__and2_1
X_09565_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ net823 net235 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout163_X net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06777_ net422 _00985_ net195 _00971_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08516_ net1079 _03979_ vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__xor2_1
X_05728_ net474 _01432_ _01431_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ net940 net202 _04624_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__o21a_1
XANTENNA__07113__A2 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ _03630_ _03906_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__o21ai_1
X_05659_ _01322_ _01326_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08378_ _00711_ _00727_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08074__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07329_ _02943_ _01040_ _00964_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10340_ clknet_leaf_25_wb_clk_i _00280_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_115_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ clknet_leaf_8_wb_clk_i _00263_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09574__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
Xfanout461 net463 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_4
Xfanout472 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\] vssd1
+ vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_2
XFILLER_0_45_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout483 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07561__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06560__B1 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06177__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05081__A _00807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10924__668 vssd1 vssd1 vccd1 vccd1 net668 _10924__668/LO sky130_fd_sc_hd__conb_1
XFILLER_0_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06863__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout90 _01606_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_2
X_10607_ clknet_leaf_35_wb_clk_i _00471_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ clknet_leaf_30_wb_clk_i _00406_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10469_ clknet_leaf_13_wb_clk_i net827 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_back
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07736__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06640__A _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09951__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_04961_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] vssd1 vssd1
+ vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
X_06700_ _01740_ _02283_ _02372_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__o21ai_1
X_07680_ net200 _01700_ _01723_ _02829_ _02835_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__o311a_1
XANTENNA__06639__X _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06631_ _02109_ _02301_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09350_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__or2_1
X_06562_ _02148_ net249 _02176_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_47_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08301_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__and2b_1
X_10825__500 vssd1 vssd1 vccd1 vccd1 _10825__500/HI net500 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_47_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05513_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _01223_ _01201_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a211o_1
X_09281_ net226 _04473_ _04474_ net396 net1158 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06493_ net130 net123 _01684_ _02061_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__o31a_1
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09398__A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\] _03710_
+ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_99_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05444_ _01023_ _01080_ _01090_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_16_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06815__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08163_ _03635_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_136_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05375_ net190 _01004_ _01014_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06534__B _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07114_ _01811_ _02282_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ _03599_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ net229 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload60 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinv_4
Xclkload71 clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__inv_8
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07045_ net282 _00757_ _02697_ _02699_ _01920_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_73_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06550__A _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07031__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__or4b_1
XANTENNA__05166__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ _03500_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__nand2_1
XANTENNA__06549__X _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _03345_ _03399_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__and3_1
X_09617_ _04688_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06829_ _02498_ _02499_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__nor2_2
XFILLER_0_35_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ net904 net203 _04653_ vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07098__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09479_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] _00667_
+ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05900__Y _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06845__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08047__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10993__633 vssd1 vssd1 vccd1 vccd1 _10993__633/HI net633 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ clknet_leaf_50_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[0\]
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10254_ clknet_leaf_4_wb_clk_i _00246_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06460__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10172__RESET_B net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10185_ clknet_leaf_78_wb_clk_i net448 net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10101__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07573__A2 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_1
Xfanout291 _03033_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08038__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05160_ _00848_ _00849_ _00854_ _00872_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09946__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05091_ net479 _00811_ _00816_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__and3_2
XFILLER_0_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08061__S net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09002__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08850_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ net293 net291 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ _04185_ vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07801_ _01049_ net99 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__xnor2_1
X_08781_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _04141_ vssd1 vssd1
+ vccd1 vccd1 _04142_ sky130_fd_sc_hd__or4_2
X_05993_ _01643_ net169 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07732_ _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__nand2b_1
X_04944_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] vssd1 vssd1 vccd1
+ vccd1 _00684_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05714__A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07663_ _03212_ _03216_ _03219_ _03220_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__or4b_1
XFILLER_0_79_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09402_ _00813_ _00815_ _02961_ _04555_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__or4_1
X_06614_ _02269_ _02284_ _02285_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__o22a_1
XANTENNA__05878__A2 _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ _03152_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09333_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06545_ net210 _01655_ _02054_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_X clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout240_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout338_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06476_ net86 _02148_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__nand2_4
XFILLER_0_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08215_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] net457
+ _01270_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__nand3b_1
XANTENNA__08029__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05427_ _01071_ _01096_ _01104_ _01070_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__o22a_1
X_09195_ net1151 net401 net206 _04411_ vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__a22o_1
X_10977__617 vssd1 vssd1 vccd1 vccd1 _10977__617/HI net617 sky130_fd_sc_hd__conb_1
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _03631_ _03632_ _03629_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05358_ _00669_ net393 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08077_ net410 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05289_ net191 _01001_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07028_ net285 _00754_ net83 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold11 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04248_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__o21ai_1
Xhold44 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\]
+ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[4\] vssd1 vssd1
+ vccd1 vccd1 net768 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc vssd1 vssd1
+ vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06439__B _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05869__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872_ net547 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05997__C _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06455__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10353__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ clknet_leaf_43_wb_clk_i net777 net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10237_ clknet_leaf_74_wb_clk_i net730 net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_10168_ clknet_leaf_26_wb_clk_i _00178_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10099_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.buttonHighlightDetect
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_63_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06330_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\] _02004_ _02005_
+ _01998_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__or4b_1
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06261_ _00684_ _01574_ _01575_ _01937_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a31o_1
XANTENNA__07482__A1 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08000_ _03550_ _03551_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__xnor2_1
X_05212_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00925_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06192_ net184 net176 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__nand2_4
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06037__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] vssd1 vssd1 vccd1
+ vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
X_05143_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07196__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ net7 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
X_05074_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1 vccd1 vccd1
+ _00802_ sky130_fd_sc_hd__or2_1
XANTENNA__05709__A _01421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08902_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] _04216_ net259
+ vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ net845 net151 net149 _04876_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a22o_1
X_08833_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] _04142_
+ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout190_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__C1 _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] net1033 net238 vssd1
+ vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
X_05976_ net197 _01667_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _00754_ _01961_ _03113_ _03270_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__o211ai_1
X_04927_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
X_08695_ net258 _01240_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__a21o_1
XANTENNA__06259__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05163__B _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ _01728_ _02154_ _01874_ net254 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_105_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07577_ net147 net168 net105 vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__and3_1
X_09316_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__inv_2
X_06528_ _01705_ _02039_ _02060_ _02102_ _02200_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04449_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06459_ _02131_ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09178_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07818__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06579__A3 _02149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07537__C _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__07528__A2 _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ clknet_leaf_33_wb_clk_i _00101_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05906__X _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05354__A _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__A3 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10924_ net668 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_0_39_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ net530 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10786_ clknet_leaf_1_wb_clk_i _00607_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10208__Q team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07216__A1 _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06019__A2 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07728__B net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05248__B _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06727__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05830_ _01520_ _01523_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05761_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\] vssd1 vssd1 vccd1
+ vccd1 _01460_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_85_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07500_ _02250_ _02673_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08480_ _03947_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2_1
X_05692_ net434 _01404_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07431_ _03013_ net230 _03012_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[17\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_18_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06366__Y _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07362_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05711__B _01423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09101_ net208 _04341_ _04343_ net397 net779 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06313_ net215 _01969_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07293_ _02923_ _02924_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ _04286_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__and3_1
X_06244_ net275 _01920_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__and2_2
XANTENNA__06382__X _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06823__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\] vssd1
+ vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold311 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] vssd1
+ vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ net186 net114 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout203_A _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold333 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08955__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold344 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_right vssd1
+ vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__dlygate4sd3_1
X_05126_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ _00838_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__and3_1
Xhold355 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold366 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\] vssd1 vssd1 vccd1
+ vccd1 net1035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold377 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold399 _00019_ vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__dlygate4sd3_1
X_05057_ _00772_ _00784_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__nor2_1
X_09934_ net1104 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input8_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ net234 _04228_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__and3_1
XANTENNA__06718__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ net192 _04165_ vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] _04815_ vssd1
+ vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or2_1
X_08747_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ net239 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__mux2_1
X_05959_ _01574_ _01575_ net144 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a21o_4
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold150_A team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ _04080_ _04102_ _04084_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06497__A2 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ _03181_ _03185_ _03186_ _02734_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ clknet_leaf_35_wb_clk_i _00504_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ clknet_leaf_11_wb_clk_i _00439_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08643__B1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08946__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05068__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ clknet_leaf_32_wb_clk_i net1023 net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05355__Y _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__A2 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10702__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10140__D team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06908__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ net572 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA__07685__A1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ net513 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__05250__C team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10769_ clknet_leaf_66_wb_clk_i _00590_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07739__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06362__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06412__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09969__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout109 _01615_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_4
X_07980_ _01679_ _03492_ _03495_ _03534_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06931_ _02543_ _02548_ _02559_ _02471_ net95 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__o32a_1
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09650_ _04713_ _04711_ net1127 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
X_06862_ _02494_ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__nand2_1
XANTENNA__06176__B2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08601_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01239_ vssd1
+ vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05813_ _01492_ _01504_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__xor2_1
X_09581_ _01793_ _03992_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nor2_2
XANTENNA__10382__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05923__A1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06793_ _02444_ _02456_ _02464_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08532_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\]
+ _03985_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\] vssd1 vssd1
+ vccd1 vccd1 _03991_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05744_ _00766_ _01444_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07676__A1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] net460
+ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__nand2_1
XANTENNA__07676__B2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05675_ _01344_ _01387_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ _02999_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ net459 _03868_ _03840_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07345_ net414 _02953_ _02954_ _00964_ _02955_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_col
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout320_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout418_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07276_ _02912_ _02913_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[13\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06553__A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09015_ net247 _04277_ _04278_ net404 net1065 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06227_ _01838_ _01902_ _01905_ _01906_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold130 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\] vssd1
+ vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06158_ _01835_ _01836_ _01838_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__or3_1
Xhold141 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold152 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[2\]
+ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__dlygate4sd3_1
X_05109_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ _00817_ _00823_ net1067 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold174 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\] vssd1 vssd1
+ vccd1 vccd1 net843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold185 _00498_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__dlygate4sd3_1
X_06089_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\] vssd1 vssd1 vccd1
+ vccd1 _01772_ sky130_fd_sc_hd__or3_1
Xhold196 team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\] vssd1 vssd1 vccd1
+ vccd1 net865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07384__A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] _01781_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\] vssd1 vssd1 vccd1
+ vccd1 _04898_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_126_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ net264 _04852_ _04853_ net243 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a32o_1
XANTENNA__10400__SET_B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09779_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] _04803_ vssd1
+ vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_122_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07831__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__B1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07323__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07667__A1 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07667__B2 _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10842__517 vssd1 vssd1 vccd1 vccd1 _10842__517/HI net517 sky130_fd_sc_hd__conb_1
XFILLER_0_14_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ clknet_leaf_38_wb_clk_i _00487_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ clknet_leaf_11_wb_clk_i _00422_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10485_ clknet_leaf_28_wb_clk_i _00353_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10255__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09041__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10135__D team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07658__A1 _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08855__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09949__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05460_ net393 _01166_ _01172_ _01162_ _01165_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05391_ net431 _00967_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07130_ _01694_ net163 _02775_ _02767_ _02762_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06373__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07061_ _01639_ _02714_ _02335_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_97_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06012_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07963_ _03398_ _03401_ _03516_ _03517_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\] _04742_ vssd1 vssd1
+ vccd1 vccd1 _04749_ sky130_fd_sc_hd__and4_1
X_06914_ _02535_ _02584_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__nand2_1
X_07894_ net106 _01692_ net183 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] _04698_ vssd1
+ vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__or2_1
X_06845_ net197 _02500_ _02515_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__o21a_1
X_09564_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ net784 net235 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
X_06776_ _00984_ net173 _02447_ net183 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08515_ _00698_ _03976_ _03979_ vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__a21oi_1
X_05727_ _01432_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
X_09495_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ net266 _04623_ net288 net218 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout156_X net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08446_ _03908_ _03919_ net489 _03753_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05658_ _01255_ _01278_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__nand2_1
X_10945__585 vssd1 vssd1 vccd1 vccd1 _10945__585/HI net585 sky130_fd_sc_hd__conb_1
XFILLER_0_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ _03835_ _03852_ net488 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05589_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] vssd1 vssd1 vccd1
+ vccd1 _01302_ sky130_fd_sc_hd__or3b_2
XFILLER_0_18_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07328_ _02942_ _02419_ _01109_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07259_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ _02900_ _02902_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10270_ clknet_leaf_7_wb_clk_i _00262_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07585__B1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[2\] vssd1 vssd1 vccd1
+ vccd1 net440 sky130_fd_sc_hd__clkbuf_2
Xfanout451 net452 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_2
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
Xfanout473 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\] vssd1
+ vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_2
Xfanout484 net486 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_2
XFILLER_0_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06458__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06560__A1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06177__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08225__A_N net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06464__Y _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout91 net92 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_2
X_10606_ clknet_leaf_35_wb_clk_i _00470_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06193__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10537_ clknet_leaf_30_wb_clk_i _00405_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_17_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ clknet_leaf_13_wb_clk_i net778 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_select
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07736__B _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06379__A1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10399_ clknet_leaf_17_wb_clk_i net673 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07591__A3 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04960_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\] vssd1 vssd1
+ vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06000__B1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ _02291_ _02299_ _02302_ _02259_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a31o_1
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06551__A1 _02220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06561_ _02067_ _02150_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08300_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05512_ net420 _01221_ _01222_ _01224_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a22o_1
X_09280_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06492_ _02076_ _02155_ _02153_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_47_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08231_ _03708_ _03709_ _03702_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__o21a_1
X_05443_ _01061_ _01070_ _01094_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_99_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06374__Y _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06815__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08162_ net466 _03639_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nand2_1
XANTENNA__08056__B2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05374_ net191 _01013_ _01086_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07113_ _01634_ _02332_ _02766_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a21oi_4
X_08093_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ _00814_ net476 vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout116_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload50 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07044_ _02088_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__nor2_2
Xclkload61 clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_8
Xclkload72 clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06831__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06550__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__or2_1
XANTENNA__05166__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ net270 _03414_ _03416_ net272 vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__o22ai_1
XANTENNA__09859__A2 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__A _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _01145_ net110 _03431_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\] _04682_ vssd1 vssd1
+ vccd1 vccd1 _04688_ sky130_fd_sc_hd__and4_1
X_06828_ net427 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1 vssd1
+ vccd1 vccd1 _02499_ sky130_fd_sc_hd__nor2_1
XANTENNA__06542__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05182__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09547_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ net268 net290 net222 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a211o_1
X_06759_ net216 _02419_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__nand2_1
X_09478_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ net218 _04605_ net886 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08429_ _03639_ _03899_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_117_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08047__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__inv_12
XFILLER_0_74_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10322_ clknet_leaf_25_wb_clk_i net738 net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_131_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10253_ clknet_leaf_4_wb_clk_i _00245_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06460__B _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05357__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ clknet_leaf_82_wb_clk_i net452 net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05033__A1 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout270 _01622_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07572__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout292 _03033_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08955__X _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10848__523 vssd1 vssd1 vccd1 vccd1 _10848__523/HI net523 sky130_fd_sc_hd__conb_1
XFILLER_0_9_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06475__X _02149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08038__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06049__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05819__X _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05090_ _00813_ _00815_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06370__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10935__584 vssd1 vssd1 vccd1 vccd1 _10935__584/HI net584 sky130_fd_sc_hd__conb_1
X_07800_ _01078_ net93 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08780_ net399 _01453_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05992_ net178 net169 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__nor2_2
XANTENNA__06772__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06772__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ _01105_ net271 _01625_ _01636_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a31o_1
X_04943_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] vssd1
+ vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XANTENNA__05980__C1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07662_ _01904_ _02765_ _03071_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__or3_1
XANTENNA__05714__B _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ _02962_ _03592_ _04556_ _02963_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__o2bb2a_1
X_06613_ _01653_ _02270_ net250 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a21o_1
XANTENNA__05878__A3 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07593_ net87 _02298_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_66_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09332_ net223 net395 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__mux2_1
X_06544_ net96 _02131_ _02215_ _02217_ _02211_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a41o_1
XFILLER_0_133_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05730__A _00711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09263_ net227 _04461_ _04462_ net403 net1168 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06475_ net86 _02148_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout233_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08214_ _01293_ _03676_ _03692_ net458 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__o22a_1
XANTENNA__10367__SET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08029__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05426_ _00966_ _01081_ _01050_ _01036_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__a2bb2o_1
X_09194_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08145_ net467 net469 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nor2_2
X_05357_ net189 _01005_ _01021_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout400_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout119_X net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08076_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ _03024_ net295 net1053 _03590_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__a221o_1
XANTENNA__06561__A _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05288_ _00996_ _01000_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07027_ _02677_ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09872__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold12 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__o21a_1
Xhold34 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _01078_ net198 _03312_ _01068_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__o22a_1
Xhold78 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi vssd1 vssd1
+ vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06515__A1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ net546 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09465__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960__600 vssd1 vssd1 vccd1 vccd1 _10960__600/HI net600 sky130_fd_sc_hd__conb_1
XFILLER_0_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09768__A1 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07567__A _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10305_ clknet_leaf_42_wb_clk_i _00043_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10236_ clknet_leaf_75_wb_clk_i net710 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10167_ clknet_leaf_55_wb_clk_i _00177_ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10098_ clknet_leaf_74_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[3\]
+ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10889__645 vssd1 vssd1 vccd1 vccd1 net645 _10889__645/LO sky130_fd_sc_hd__conb_1
XFILLER_0_107_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07703__B1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06260_ _01677_ _01936_ net456 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07482__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05211_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00924_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_133_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06191_ net215 net101 net92 net197 _01871_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05142_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__nand2_1
Xhold504 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08072__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06381__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07196__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09950_ net461 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
X_05073_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1 vccd1 vccd1
+ _00801_ sky130_fd_sc_hd__nand2_1
X_08901_ _01404_ _04198_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09881_ _01773_ _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08832_ _04142_ _04175_ net193 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07942__B1 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05725__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
X_05975_ net256 net170 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_68_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout183_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07714_ net95 _02217_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__or2_1
X_04926_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] vssd1
+ vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
X_08694_ _04112_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07645_ _03180_ _03187_ _03191_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_105_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout448_A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ net142 net166 net162 net137 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09315_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__and3_1
X_06527_ net136 _01698_ _02056_ _02091_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout236_X net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09246_ net228 _04448_ _04450_ net406 net890 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__a32o_1
X_06458_ net201 _02112_ _02113_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__or3_1
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05409_ _01083_ _01087_ _01093_ _01098_ _01082_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__o2111a_1
X_09177_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04396_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__and2_1
XANTENNA__06681__B1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06389_ _02060_ _02061_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08128_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08059_ net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ net389 net293 vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_102_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout96_A _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
X_10021_ clknet_leaf_33_wb_clk_i _00100_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_129_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05922__X _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07850__A _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ net667 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_86_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07161__A1 _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05172__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__A3 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10854_ net529 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10785_ clknet_leaf_66_wb_clk_i _00606_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.audio
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06672__B1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06019__A3 _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10224__Q team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10219_ clknet_leaf_82_wb_clk_i _00223_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07924__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05760_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _01458_
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__or4b_1
XANTENNA__09677__A0 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05691_ net487 _00796_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__nand2_1
XANTENNA__07152__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07430_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ _03009_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06376__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07361_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09100_ _04342_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__inv_2
X_06312_ net196 _01966_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07455__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07292_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06663__X _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09031_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ _04286_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06243_ net278 net272 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__nor2_1
XANTENNA__07928__A1_N _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06174_ net210 net97 net94 net194 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
Xhold301 _00022_ vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold312 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold323 _00028_ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10244__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold334 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__dlygate4sd3_1
X_05125_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__nand2_1
XANTENNA__08955__A2 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_right vssd1
+ vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold367 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\] vssd1 vssd1 vccd1
+ vccd1 net1036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] vssd1 vssd1
+ vccd1 vccd1 net1047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\] vssd1 vssd1 vccd1
+ vccd1 net1058 sky130_fd_sc_hd__dlygate4sd3_1
X_05056_ net1030 _00774_ _00784_ _00786_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[5\]
+ sky130_fd_sc_hd__o31ai_1
X_09933_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ net825 net258 _04864_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__a21o_1
XANTENNA__06718__A1 _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ net972 _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_107_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _04811_ _04814_ _04816_ _04808_ net1167 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_29_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08746_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ net239 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__mux2_1
X_05958_ net144 net133 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_124_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04909_ net277 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XANTENNA__07143__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05889_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] _01579_
+ _01581_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__and3_2
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _04089_ _04092_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07628_ _01660_ _02061_ _03183_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__a21bo_1
XANTENNA__05902__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ _02135_ _02140_ _02150_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__a21oi_2
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10570_ clknet_leaf_9_wb_clk_i _00438_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09229_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04435_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08946__A2 _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout99_X net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06709__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__B2 _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ clknet_leaf_32_wb_clk_i _00024_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05067__D_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06908__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10906_ net571 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XANTENNA__07685__A2 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06196__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ net512 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_7_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10768_ clknet_leaf_59_wb_clk_i _00589_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10699_ clknet_leaf_66_wb_clk_i _00530_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06362__C _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05259__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06930_ _02533_ _02585_ _02600_ _02569_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06861_ _02530_ _02531_ _02475_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06176__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03623_ net751 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__o21a_1
X_05812_ _01492_ _01504_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__xnor2_1
X_09580_ _01793_ _03967_ _03976_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__o21ai_2
X_06792_ net113 _02458_ _02463_ _02457_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05923__A2 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\] _03985_ vssd1 vssd1
+ vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand4_1
X_05743_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ _00775_ _00652_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07852__A1_N net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08462_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] _03686_
+ _03688_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__a21oi_1
X_05674_ net417 _01258_ _01381_ _01386_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__a211o_1
XANTENNA__07676__A2 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07413_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ _02998_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\] vssd1
+ vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__a31o_1
X_08393_ _01257_ _03728_ _03867_ net460 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_86_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout146_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07489__X _03050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07344_ net491 net414 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07275_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout313_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09014_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__or2_1
X_06226_ net97 _01878_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08389__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06157_ net95 _01831_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__nor2_1
Xhold120 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[8\] vssd1 vssd1
+ vccd1 vccd1 net789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold142 net54 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold153 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__dlygate4sd3_1
X_05108_ net1024 _00817_ _00823_ net1038 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__a22o_1
Xhold164 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\] vssd1 vssd1
+ vccd1 vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\] vssd1 vssd1
+ vccd1 vccd1 net844 sky130_fd_sc_hd__dlygate4sd3_1
X_06088_ _00654_ _01771_ _01411_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21oi_1
Xhold186 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] vssd1 vssd1
+ vccd1 vccd1 net855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ net1097 net152 net150 _04897_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05039_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__nand4_1
XANTENNA__07384__B _01475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04850_ vssd1
+ vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09778_ _04799_ _04800_ _04801_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_122_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08729_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__mux2_1
XANTENNA__07116__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10881__556 vssd1 vssd1 vccd1 vccd1 _10881__556/HI net556 sky130_fd_sc_hd__conb_1
X_10622_ clknet_leaf_38_wb_clk_i _00486_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10166__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ clknet_leaf_12_wb_clk_i _00421_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10484_ clknet_leaf_26_wb_clk_i _00352_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input31_X net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__X _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05823__A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07107__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07107__B2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07658__A2 _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05390_ net189 _01013_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_31_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07060_ _01639_ _02713_ _02714_ _02686_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_97_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06011_ net126 _01683_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__A _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07043__B1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07962_ net257 _01621_ _03392_ _03427_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_71_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\] _04745_ vssd1
+ vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__nor2_1
X_06913_ _00751_ _02486_ _02539_ _02537_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06149__A2 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ _03306_ _03446_ _03447_ _03445_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__or4b_1
X_09632_ net1090 _04698_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__nor2_1
X_06844_ net211 _02511_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09563_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ net831 net241 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
X_06775_ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout263_A _00746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] _00657_ _01793_
+ _03977_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a31o_1
X_05726_ _01108_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back vssd1
+ vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__or3b_2
X_09494_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ _00667_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06267__C net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08445_ net462 _03713_ _03918_ _03911_ net411 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a311o_1
X_05657_ _01278_ _01369_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08376_ net485 _03846_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__or3_1
X_05588_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07327_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\] team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__mux2_1
XANTENNA__08074__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07258_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06209_ net91 _01800_ _01824_ net101 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a22o_1
X_07189_ _01717_ _01737_ _01828_ _01662_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a211o_1
XANTENNA__05908__A _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__A1 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[0\] vssd1 vssd1 vccd1
+ vccd1 net430 sky130_fd_sc_hd__buf_4
Xfanout441 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1 vccd1
+ vccd1 net441 sky130_fd_sc_hd__buf_2
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_2
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_4
Xfanout474 net483 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08938__B _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_1
XANTENNA__10322__Q team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05914__Y _01608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06739__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07334__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06560__A2 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024__643 vssd1 vssd1 vccd1 vccd1 _11024__643/HI net643 sky130_fd_sc_hd__conb_1
XFILLER_0_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout81 _02731_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_4
XFILLER_0_52_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10605_ clknet_leaf_35_wb_clk_i _00469_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout92 _01606_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10536_ clknet_leaf_30_wb_clk_i _00404_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10372__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ clknet_leaf_29_wb_clk_i net729 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_right
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06480__Y _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__B net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06379__A2 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ clknet_leaf_17_wb_clk_i net718 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07576__B2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11019_ net642 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_0_95_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06000__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06001__X _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06368__B _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05272__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ _01739_ net164 _02092_ _02155_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05511_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ _01198_ _01203_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06491_ net275 net279 _00747_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _00683_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__nand2_2
X_05442_ _01038_ _01079_ _01067_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08161_ net473 _03634_ _03639_ net466 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a31o_1
X_05373_ _01085_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
X_10905__570 vssd1 vssd1 vccd1 vccd1 _10905__570/HI net570 sky130_fd_sc_hd__conb_1
XFILLER_0_67_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07112_ _02332_ net81 _02735_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a21oi_1
X_08092_ net949 net229 _03595_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07043_ _01675_ _01828_ net199 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a21oi_1
Xclkload40 clknet_leaf_57_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_4
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload51 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__clkinv_8
Xclkload62 clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_6
XFILLER_0_113_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload73 clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_4
XANTENNA_fanout109_A _01615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06550__C _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04260_ _04262_ _04258_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__o31a_1
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ _03480_ _03486_ _03493_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a22o_1
XANTENNA__10327__SET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout380_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A3 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__B _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ _00970_ net119 net110 _01145_ _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09615_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\]
+ _04682_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 _04687_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06827_ net427 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1 vssd1
+ vccd1 vccd1 _02498_ sky130_fd_sc_hd__and2_1
XANTENNA__06542__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ net911 net204 _04652_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06758_ _02428_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05709_ _01421_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
X_09477_ net886 net203 _04611_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__o21a_1
X_06689_ net99 net90 net86 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08428_ _03662_ _03891_ _00703_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_22_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08359_ team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel _03719_ _03834_
+ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10321_ clknet_leaf_24_wb_clk_i net788 net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07329__S _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10252_ clknet_leaf_46_wb_clk_i _00244_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07558__A1 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10183_ clknet_leaf_23_wb_clk_i _00193_ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout81_X net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input39_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 _00756_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_4
Xfanout271 _01620_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_4
Xfanout282 net284 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07572__B net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10887__562 vssd1 vssd1 vccd1 vccd1 _10887__562/HI net562 sky130_fd_sc_hd__conb_1
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10110__RESET_B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07494__B1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06049__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10519_ clknet_leaf_29_wb_clk_i _00387_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08746__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05991_ net210 net179 _01663_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a21o_2
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07730_ net108 _03280_ _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__or3b_2
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04942_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\] vssd1 vssd1
+ vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XANTENNA__05980__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07661_ _02829_ _03213_ _03218_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_49_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05714__C _01423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ _02959_ _02961_ _02964_ team_07_WB.instance_to_wrap.ssdec_ss _04556_ vssd1
+ vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__a221o_1
X_06612_ _01720_ _02021_ _02271_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ _01664_ _01669_ _03149_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09331_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ net6 net322 _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06543_ net89 _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09262_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ _04459_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06474_ _01596_ _01603_ _01598_ _01590_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__o211a_4
XFILLER_0_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ _01281_ _03679_ _03691_ net459 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_62_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05425_ net432 _01099_ _01113_ _01085_ _01137_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__a221o_1
X_09193_ net206 _04409_ _04410_ net401 net1162 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07497__X _03057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nand2_2
X_05356_ _00967_ _01062_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__or2_1
XANTENNA__08434__C1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__A1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08075_ net454 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__and2b_1
X_05287_ _00675_ _00999_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_112_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06561__B _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07026_ _02678_ _02680_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] net820
+ net445 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
Xhold24 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
X_10914__658 vssd1 vssd1 vccd1 vccd1 net658 _10914__658/LO sky130_fd_sc_hd__conb_1
Xhold35 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07928_ _01068_ _03312_ net187 _01091_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a2bb2o_1
Xhold57 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\] vssd1 vssd1
+ vccd1 vccd1 net737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07859_ _03299_ _03413_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__or2_1
XANTENNA__05318__A3 _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ net545 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ net267 _04643_ net289 net220 vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06279__A1 _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07491__A3 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07567__B _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06451__A1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ clknet_leaf_24_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[17\]
+ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06451__B2 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10235_ clknet_leaf_74_wb_clk_i net712 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10709__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06203__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06203__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10166_ clknet_leaf_58_wb_clk_i _00176_ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_10097_ clknet_leaf_74_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[2\]
+ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10362__RESET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07703__B2 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05390__X _01103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10999_ net636 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_44_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07467__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05210_ _00919_ _00920_ _00921_ _00922_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_133_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06190_ net186 net114 _01866_ _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_72_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06662__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05141_ _00850_ _00851_ _00852_ _00853_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold505 team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\] vssd1 vssd1 vccd1
+ vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05072_ net423 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1 vssd1
+ vccd1 vccd1 _00800_ sky130_fd_sc_hd__xor2_1
XANTENNA__07196__C _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08900_ _04215_ net924 _04209_ vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09880_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] _01772_ vssd1
+ vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nand2_1
XANTENNA__10090__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08831_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\]
+ _04141_ net877 vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09931__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__A1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__B2 _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
X_05974_ net179 net177 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__or2_2
X_07713_ _03256_ _03258_ _03268_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_68_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04925_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] vssd1
+ vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
X_08693_ net242 _04113_ _04040_ _01759_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout176_A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10983__623 vssd1 vssd1 vccd1 vccd1 _10983__623/HI net623 sky130_fd_sc_hd__conb_1
X_07644_ _03074_ _03192_ _03195_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_105_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06837__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07575_ _01686_ _02263_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout343_A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ _04491_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06526_ _01687_ _01690_ _02047_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09245_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__inv_2
X_06457_ _01711_ _02089_ _02050_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05408_ _01111_ _01112_ _01119_ _01120_ _01073_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__o2111a_1
X_09176_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04396_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__or2_1
X_06388_ _02061_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__inv_2
XANTENNA__08958__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08127_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\] _03613_
+ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05339_ net190 _01004_ _01005_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__nor3_2
XFILLER_0_32_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08058_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net291 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07009_ _02661_ _02665_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__and2_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
X_10020_ clknet_leaf_33_wb_clk_i net950 net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout89_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ net666 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XANTENNA__07850__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05172__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10853_ net528 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_39_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08646__C1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ clknet_leaf_64_wb_clk_i _00605_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10218_ clknet_leaf_79_wb_clk_i _00222_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05545__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ clknet_leaf_17_wb_clk_i net705 net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_10967__607 vssd1 vssd1 vccd1 vccd1 _10967__607/HI net607 sky130_fd_sc_hd__conb_1
XANTENNA__09126__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05690_ net487 _00796_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07360_ _02968_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_fl_enable
+ sky130_fd_sc_hd__inv_2
XFILLER_0_128_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06311_ net196 _01966_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06521__A2_N _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07291_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ _02922_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09030_ net248 _04288_ _04289_ net404 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__a32o_1
X_06242_ _01827_ _01847_ _01918_ _01919_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[3\]
+ sky130_fd_sc_hd__and4_1
XANTENNA__06392__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06173_ net211 net95 _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold302 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\] vssd1 vssd1
+ vccd1 vccd1 net971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\] vssd1 vssd1 vccd1
+ vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05124_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ _00835_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__a21o_1
Xhold324 net52 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold346 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] vssd1 vssd1
+ vccd1 vccd1 net1015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\] vssd1 vssd1 vccd1
+ vccd1 net1026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\] vssd1 vssd1 vccd1
+ vccd1 net1037 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net408 _01787_ net843 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__o21a_1
X_05055_ _00766_ _00774_ _00785_ net1030 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold379 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] vssd1 vssd1
+ vccd1 vccd1 net1048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09863_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ net234 _04228_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__and3_1
XANTENNA__06179__B1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__RESET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08814_ _04163_ _04164_ net192 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__a21oi_1
X_09794_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ net239 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
X_05957_ net130 net124 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_124_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04908_ net284 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
X_08676_ _04099_ _04101_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__a21o_1
X_05888_ _01578_ _01580_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07627_ _02171_ _03184_ _03183_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07558_ _01921_ _02214_ _01618_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06509_ _00750_ _01611_ _02042_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07489_ _01730_ _02082_ _03048_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__o211a_1
XANTENNA__08643__A2 _01475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09228_ net228 _04436_ _04437_ net406 net917 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09159_ net206 _04385_ _04386_ net402 net857 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08946__A3 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05917__Y _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06709__A2 _02149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ clknet_leaf_36_wb_clk_i _00023_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input21_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07861__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06477__A _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05381__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10905_ net570 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10836_ net511 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ clknet_leaf_59_wb_clk_i _00588_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06645__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06645__B2 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10698_ clknet_leaf_65_wb_clk_i _00529_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07755__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06860_ net92 _02474_ _02529_ _01615_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_52_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08867__A team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05811_ _00713_ _01492_ net215 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__or3_1
X_06791_ net113 _02458_ _02462_ net120 _02461_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__o221a_1
X_08530_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\] _03978_ vssd1
+ vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05742_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] _00775_ _00783_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\] vssd1 vssd1 vccd1 vccd1
+ _01443_ sky130_fd_sc_hd__a31o_1
XANTENNA__08322__A1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08461_ net806 net129 _03933_ vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05673_ _01276_ _01279_ _01300_ _01385_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__a31o_1
X_07412_ net978 _02999_ _03001_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[10\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07450__A_N net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07343_ _01109_ _02953_ _00710_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_34_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06393__Y _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09210__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ _01389_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__nand2_1
X_06225_ _01812_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout306_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold110 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ net91 _01834_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__nand2_1
Xhold121 _00135_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold143 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__dlygate4sd3_1
X_05107_ net475 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ _00821_ _00817_ net968 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a32o_1
XANTENNA__07061__A1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold176 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] vssd1 vssd1
+ vccd1 vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
X_06087_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] _01771_ _01411_
+ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21o_1
Xhold187 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] vssd1 vssd1
+ vccd1 vccd1 net856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] _01781_
+ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__xnor2_1
X_05038_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__and4b_1
XFILLER_0_10_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09846_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04850_ vssd1
+ vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07681__A _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__or4bb_1
XANTENNA__06572__B1 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\]
+ _02651_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] vssd1
+ vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ net1094 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05913__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07116__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08659_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ _04049_ _04051_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__o22a_1
XANTENNA__06324__B1 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06584__X team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10621_ clknet_leaf_38_wb_clk_i _00485_ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10771__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ clknet_leaf_11_wb_clk_i _00420_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10483_ clknet_leaf_28_wb_clk_i _00351_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07052__A1 _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10135__RESET_B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input24_X net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06563__B1 _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05382__Y _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05823__B _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08855__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06866__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08068__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ net494 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06618__A1 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06618__B2 _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06010_ net134 _01685_ net142 _01683_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07043__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__B _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07961_ _01689_ _03380_ _03388_ _01679_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09700_ _04734_ _04746_ _04747_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06912_ _01650_ _02493_ _02575_ _02582_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__or4_1
X_07892_ _01091_ net172 vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__xor2_1
X_09631_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ _04696_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06843_ net197 _02500_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__nor2_1
X_09562_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ net809 net241 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06774_ net421 _00973_ _00985_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__o21a_1
X_08513_ _00698_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05725_ net474 net490 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__nor2_1
X_09493_ net916 net203 _04622_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__o21a_1
XANTENNA__09766__B1_N _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08444_ net484 _03881_ _03917_ _03722_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_33_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05656_ _01280_ _01331_ _01337_ _01342_ _01368_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__a41o_1
XFILLER_0_72_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ _03709_ _03848_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05587_ _01295_ _01299_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07326_ _02939_ _02941_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[1\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07257_ _02898_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ _02901_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06208_ _01837_ _01845_ _01835_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07188_ _02277_ _02836_ _02829_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06139_ _01809_ _01817_ _01818_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a31o_1
XANTENNA__07346__A_N _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__A2 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout420 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\] vssd1
+ vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout431 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[2\] vssd1 vssd1
+ vccd1 vccd1 net431 sky130_fd_sc_hd__buf_4
XFILLER_0_100_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout442 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[0\] vssd1 vssd1 vccd1
+ vccd1 net442 sky130_fd_sc_hd__buf_2
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_2
Xfanout464 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.frameBufferLowNibble
+ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_8
Xfanout475 net476 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05924__A _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout486 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
X_09829_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] _04838_ vssd1
+ vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__and2_1
XANTENNA__06545__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08300__A _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06739__B net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08298__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05520__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10604_ clknet_leaf_35_wb_clk_i _00468_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout82 _02731_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_2
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_4
XFILLER_0_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10535_ clknet_leaf_30_wb_clk_i _00403_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10466_ clknet_leaf_29_wb_clk_i net719 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_left
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06490__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07025__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10397_ clknet_leaf_17_wb_clk_i net876 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06379__A3 _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11018_ net386 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_26_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06000__A2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08864__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05510_ net420 net419 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__nand2b_4
X_06490_ net282 net274 _00748_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__and3_2
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05441_ _01030_ _01097_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ net469 _03644_ _03634_ vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__mux2_1
X_05372_ net189 _01014_ _01019_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__nor3_2
XFILLER_0_16_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07111_ _02764_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ _03598_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ net229 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload30 clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_6
XFILLER_0_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload41 clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__inv_6
X_07042_ _02086_ _02696_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload52 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__clkinv_4
Xclkload63 clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__inv_8
XFILLER_0_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload74 clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload74/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_73_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08993_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04261_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832__507 vssd1 vssd1 vccd1 vccd1 _10832__507/HI net507 sky130_fd_sc_hd__conb_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07944_ _03496_ _03498_ _03495_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10951__591 vssd1 vssd1 vccd1 vccd1 _10951__591/HI net591 sky130_fd_sc_hd__conb_1
X_07875_ _00970_ net119 _03349_ _03423_ _03348_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09614_ _04685_ _04686_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__nand2_1
X_06826_ _02495_ _02496_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09545_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ net268 net290 net222 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06757_ net252 _02427_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout161_X net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05708_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _01419_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__or3_2
X_09476_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ net266 net287 net218 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a211o_1
XANTENNA__06575__A _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06688_ _01223_ _01413_ _02324_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a21oi_1
X_08427_ _03657_ _03755_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__or3b_1
X_05639_ _01350_ _01351_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08358_ net486 net412 _03719_ _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload2 clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_22_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07309_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ _03632_ _03661_ _03765_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ clknet_leaf_24_wb_clk_i net826 net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10251_ clknet_leaf_74_wb_clk_i _00243_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05357__C _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ clknet_leaf_23_wb_clk_i _00192_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout250 net251 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_4
Xfanout261 _00756_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 _00752_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_4
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07572__C net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09560__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07494__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06049__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10518_ clknet_leaf_29_wb_clk_i _00386_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08205__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10449_ clknet_leaf_24_wb_clk_i _00333_ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_90_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05990_ net210 net179 _01663_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a21oi_4
X_04941_ net437 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07660_ net130 _01676_ net165 _02835_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_49_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07182__B1 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06611_ _02013_ _02073_ _02276_ _02282_ net250 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a221oi_4
X_07591_ _01543_ net143 _01658_ _03077_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__o31ai_1
X_09330_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ net6 _04312_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a21oi_1
X_06542_ net119 net271 net112 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_66_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06395__A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04908__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ _04459_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06473_ _02143_ _02145_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_138_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08212_ net460 _03689_ _03690_ _01283_ _03681_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__o32a_1
X_05424_ _01030_ _01048_ _01056_ _01034_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__a2bb2o_1
X_09192_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ _04407_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ _00702_ _03628_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__or2_2
XFILLER_0_71_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05355_ net296 _01067_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__nor2_4
XFILLER_0_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout121_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__A2 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ net392 net295 net1033 _03589_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__a221o_1
X_05286_ _00976_ _00997_ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07025_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] net298 net394 _02679_
+ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold14 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] net835
+ net445 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
Xhold25 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05474__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold47 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\] vssd1 vssd1
+ vccd1 vccd1 net727 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ net296 _01665_ _03310_ _03481_ _03303_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__o32a_1
Xhold69 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06289__B net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07858_ net276 _03292_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__nand2_1
XANTENNA__07173__B1 _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ _02479_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__inv_2
X_07789_ _01050_ _01590_ _01598_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06576__Y _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09528_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] _00666_
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] vssd1 vssd1
+ vccd1 vccd1 _04643_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09459_ net927 net202 _04601_ _04602_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__o22a_1
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07228__A1 _02081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07228__B2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08025__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05001__X _00738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10303_ clknet_leaf_25_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[16\]
+ net357 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10234_ clknet_leaf_71_wb_clk_i net692 net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_10165_ clknet_leaf_20_wb_clk_i _00175_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05384__A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ clknet_leaf_74_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\]
+ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07164__B1 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10998_ net387 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_44_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07467__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07758__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06662__B _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05140_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] vssd1 vssd1
+ vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05071_ _00672_ net429 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_41_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08830_ _04173_ _04174_ net193 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07942__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08761_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__mux2_1
XANTENNA__10385__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05973_ net181 net174 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__nor2_1
X_07712_ _03260_ _03264_ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__and3_2
X_04924_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08692_ _01243_ _01251_ _04035_ _01250_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__o211a_1
XANTENNA__07155__B1 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07643_ _01730_ _02765_ _03073_ _03105_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__o32a_1
XFILLER_0_79_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06902__B1 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07574_ _02033_ _02040_ net162 _02836_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_24_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09313_ net225 _04496_ _04497_ net401 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a32o_1
X_06525_ _02139_ _02195_ _02196_ _02198_ _02193_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a311o_1
XFILLER_0_8_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09244_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06456_ _02059_ _02072_ _02093_ _02128_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__o31a_1
XFILLER_0_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05407_ _01106_ _01107_ _01115_ _01060_ _01118_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09175_ net207 _04395_ _04397_ net401 net999 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06387_ net214 net173 net137 _01684_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a31o_2
XFILLER_0_32_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08958__A1 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__or2_1
X_05338_ net393 _01049_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08057_ _03582_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net294 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10838__513 vssd1 vssd1 vccd1 vccd1 _10838__513/HI net513 sky130_fd_sc_hd__conb_1
X_05269_ net422 _00979_ net421 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07008_ _02658_ _02667_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__xor2_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08959_ _04247_ net419 _04245_ vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05932__A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ net665 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__07697__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10852_ net527 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_128_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ clknet_leaf_64_wb_clk_i _00604_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10895__651 vssd1 vssd1 vccd1 vccd1 net651 _10895__651/LO sky130_fd_sc_hd__conb_1
XFILLER_0_132_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07594__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ clknet_leaf_82_wb_clk_i _00221_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10148_ clknet_leaf_16_wb_clk_i net753 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06497__X _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ clknet_leaf_45_wb_clk_i _00137_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07152__A3 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06310_ net437 net184 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07290_ _02921_ _02922_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[6\]
+ sky130_fd_sc_hd__or2_1
XANTENNA__06112__A1 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06673__A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06241_ _01672_ _01915_ _01917_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06392__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05289__A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06172_ net210 net95 _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold303 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\] vssd1 vssd1
+ vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold314 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] vssd1 vssd1
+ vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
X_05123_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] _00833_ vssd1 vssd1
+ vccd1 vccd1 _00836_ sky130_fd_sc_hd__nand2_1
Xhold325 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\]
+ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07612__A1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold336 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\] vssd1
+ vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold347 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] vssd1 vssd1
+ vccd1 vccd1 net1016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold358 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_down vssd1
+ vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\] vssd1
+ vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net843 net333 _01788_ _04905_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__a31o_1
X_05054_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00780_ _00766_
+ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05295__Y _01008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09862_ _00726_ _03992_ _04804_ _04863_ _04861_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a41o_1
XANTENNA__06179__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06179__B2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\]
+ _04160_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__or3_1
X_09793_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_107_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] net1108 net240 vssd1
+ vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__mux2_1
X_05956_ net134 net127 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04907_ net285 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _04075_ _04100_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__a21o_1
X_05887_ _00715_ _01575_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout453_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07626_ _02786_ _03169_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07557_ _01880_ _02743_ _03113_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06508_ net98 _02180_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07488_ net134 net141 _01729_ _01743_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09227_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04430_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__a21o_1
X_06439_ _01708_ _01732_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05199__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09158_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04379_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ net903 _02672_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__xor2_1
X_09089_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04328_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07603__B2 _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ clknet_leaf_32_wb_clk_i net970 net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10904_ net569 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10835_ net510 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10766_ clknet_leaf_66_wb_clk_i _00587_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10697_ clknet_leaf_65_wb_clk_i _00528_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06004__Y _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05810_ _01494_ _01499_ _01500_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o31a_2
X_06790_ _02410_ _02415_ _02460_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__and3_1
X_05741_ _00774_ _00783_ _01442_ _00766_ net1171 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[4\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__06020__X _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08460_ _03753_ _03932_ _03927_ net129 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__o211a_1
X_05672_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] _01260_
+ _01379_ _01380_ _01383_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06333__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07411_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] _02999_
+ net477 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__o21ai_1
X_08391_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _01259_ _01284_
+ _01305_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a41o_1
XFILLER_0_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07342_ net474 net488 _00797_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07273_ _01389_ _02911_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[12\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09012_ net247 _04275_ _04276_ net404 net880 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06224_ net200 _01829_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__or2_2
XFILLER_0_60_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06155_ net91 _01834_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout201_A _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[3\] vssd1 vssd1
+ vccd1 vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold133 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__dlygate4sd3_1
X_05106_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\]
+ _00817_ _00823_ net969 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold144 _00167_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
X_06086_ _01768_ _01769_ _01770_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__or3_1
Xhold155 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[14\]
+ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[24\]
+ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ net856 net153 net149 _04896_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05037_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07962__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _04850_ _04851_ net1109 _04824_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout191_X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07681__B _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__nand4b_1
XANTENNA__06572__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06988_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _02651_
+ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__nand2_1
XANTENNA__06578__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08727_ net1011 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05939_ _01628_ _01632_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nor2_4
X_08658_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04046_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07609_ _02254_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08589_ _03606_ _04028_ net140 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10620_ clknet_leaf_38_wb_clk_i net869 net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06088__B1 _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ clknet_leaf_12_wb_clk_i _00419_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10482_ clknet_leaf_28_wb_clk_i _00350_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06260__A0 _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09563__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07760__B1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06866__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10818_ net493 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_83_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10749_ clknet_leaf_64_wb_clk_i _00579_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09568__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05838__Y _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07043__A2 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07960_ _01092_ net118 _03507_ _03508_ _03514_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_71_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06911_ _02497_ _02521_ _02578_ _02581_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_71_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07891_ net257 _03316_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__or2_1
X_09630_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\] _04696_ net1089
+ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a21oi_1
X_06842_ net197 _02500_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06554__A1 _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06554__B2 _02149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06773_ net423 net154 _01720_ _00672_ _01736_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__o221a_1
X_09561_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ net771 net241 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05724_ net1085 _00824_ _00825_ net1067 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a22o_1
X_08512_ _01793_ _03974_ _03966_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09492_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ net268 _04614_ _04621_ net222 vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a221o_1
XANTENNA__07503__B1 _03050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08700__C1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ _03738_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__nor2_1
X_05655_ _01364_ _01367_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08059__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ net487 _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09256__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__B2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05586_ _01292_ _01294_ _01296_ _01298_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07325_ _02940_ _00974_ _00964_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07256_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06207_ _01887_ _01847_ _01827_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[0\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_115_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07187_ _02065_ net82 _02736_ _02831_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a22o_1
X_06138_ _01810_ _01814_ _01816_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11017__641 vssd1 vssd1 vccd1 vccd1 _11017__641/HI net641 sky130_fd_sc_hd__conb_1
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06069_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08073__A_N net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout421 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[2\] vssd1 vssd1
+ vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_2
Xfanout443 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[0\] vssd1 vssd1 vccd1
+ vccd1 net443 sky130_fd_sc_hd__clkbuf_2
Xfanout454 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
Xfanout465 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] vssd1
+ vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_2
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ net1031 _04836_ _04839_ _04824_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__o22a_1
Xfanout487 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_2
XANTENNA__06545__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ net244 _04786_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05940__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10603_ clknet_leaf_35_wb_clk_i net938 net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout83 _02375_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_2
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout94 _01605_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07867__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09558__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10534_ clknet_leaf_31_wb_clk_i _00402_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06481__B1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ clknet_leaf_15_wb_clk_i net732 net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_down
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06490__B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10396_ clknet_leaf_17_wb_clk_i net696 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_92_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09722__A1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ net641 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_56_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06946__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__C _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07113__Y _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05440_ _00964_ _01152_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05371_ net433 _00668_ _01067_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_56_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ _02033_ _02069_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05849__X _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08090_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ _00814_ net476 vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__o21a_1
XANTENNA__07264__A2 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload20 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_12
XFILLER_0_31_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07041_ net154 _01700_ _01828_ net199 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload31 clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload42 clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_8
XFILLER_0_70_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload53 clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_8
Xclkload64 clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__inv_8
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05297__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload75 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10026__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08992_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07972__B1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871__546 vssd1 vssd1 vccd1 vccd1 _10871__546/HI net546 sky130_fd_sc_hd__conb_1
X_07943_ _01068_ net158 _03309_ _03497_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_103_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06399__Y _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07874_ _01051_ net118 net110 _01077_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09613_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] _04664_ _04684_
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__or3_1
X_06825_ net427 net144 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09544_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ net222 _04605_ net895 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06756_ net252 _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05707_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nor2_1
X_09475_ net935 net203 _04610_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__o21a_1
X_06687_ _02354_ _02358_ _02359_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout154_X net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06575__B _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08426_ _03661_ net470 net465 vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__mux2_1
X_05638_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] vssd1 vssd1 vccd1
+ vccd1 _01351_ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08437__D1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel team_07_WB.instance_to_wrap.team_07.flagPixel
+ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__or2_1
X_05569_ net416 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01282_ sky130_fd_sc_hd__or3b_2
XFILLER_0_117_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload3 clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__inv_6
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07308_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02930_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06591__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ _00717_ net470 vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05266__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06463__B1 _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ net126 net141 _02877_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ clknet_leaf_74_wb_clk_i _00242_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10181_ clknet_leaf_20_wb_clk_i _00191_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06766__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05935__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout251 _01489_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_4
Xfanout262 _00747_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_4
Xfanout273 _00651_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
Xfanout284 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\] vssd1
+ vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_4
Xfanout295 _03026_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07494__A2 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10517_ clknet_leaf_29_wb_clk_i _00385_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05829__B _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08205__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10448_ clknet_leaf_24_wb_clk_i _00332_ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06006__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05548__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10379_ clknet_leaf_4_wb_clk_i net691 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_04940_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1 vccd1
+ vccd1 _00680_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06012__Y _01705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05980__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05717__C1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06610_ net250 _02275_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__or2_1
X_07590_ net87 _02109_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__nand2_1
XANTENNA__06676__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06541_ _01616_ _02213_ _02214_ _01618_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06395__B _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09260_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ net403 net227 _04460_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a22o_1
X_06472_ _02139_ _02141_ _02078_ _02095_ _02118_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_75_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08211_ _01285_ _03684_ _03688_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__nor3_1
X_05423_ _01131_ _01133_ _01135_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__or3_1
X_09191_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ _04407_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08142_ _00702_ _03628_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__nor2_1
X_05354_ _00966_ _01048_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__or2_4
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08073_ net454 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__and2b_1
XANTENNA__10207__RESET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05285_ _00976_ _00997_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout114_A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07024_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ net447 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08975_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] net847
+ net445 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
Xhold15 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07018__Y _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07926_ _01084_ _01652_ _01700_ _03325_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__o211ai_1
Xhold48 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07857_ _03410_ _03411_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06808_ net279 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1
+ vccd1 vccd1 _02479_ sky130_fd_sc_hd__nand2_1
XANTENNA__06586__A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07788_ _01590_ _01598_ _01050_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_27_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09527_ net936 net205 _04642_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__o21a_1
X_06739_ net425 net426 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09458_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ net265 net217 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09870__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ _03810_ _03883_ net488 vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09389_ _01415_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07228__A2 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08025__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10302_ clknet_leaf_24_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[15\]
+ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06451__A3 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958__598 vssd1 vssd1 vccd1 vccd1 _10958__598/HI net598 sky130_fd_sc_hd__conb_1
X_10233_ clknet_leaf_71_wb_clk_i net689 net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[3\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05936__Y _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ clknet_leaf_19_wb_clk_i _00174_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05411__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10095_ clknet_leaf_74_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[0\]
+ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07164__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06496__A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10997_ net387 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07120__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06007__Y _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold507 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
X_05070_ net258 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ sky130_fd_sc_hd__inv_2
XFILLER_0_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08760_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] net1177 net238 vssd1
+ vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__mux2_1
X_05972_ net253 net175 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_81_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08886__A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ _02194_ _02219_ _02738_ _03044_ _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04923_ net2 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08691_ _01749_ _01755_ _04059_ _04111_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_10_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07155__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07642_ _01737_ _02261_ _03197_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o211a_1
XANTENNA__06902__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07573_ net137 _01688_ net166 _03131_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_24_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nand2_1
X_06524_ net260 net87 _01711_ _02047_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09243_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04444_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a21o_1
XANTENNA__06666__B1 _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06455_ net263 _02030_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__or2_2
XFILLER_0_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout329_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05406_ _01071_ _01103_ _01104_ _01075_ _01076_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__o32a_1
XFILLER_0_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09174_ _04396_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__inv_2
X_06386_ _01680_ net164 _02057_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_17_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07030__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__A2 _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05337_ _00967_ _01048_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__nor2_2
X_08125_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\] _03611_
+ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or3_1
X_10920__664 vssd1 vssd1 vccd1 vccd1 net664 _10920__664/LO sky130_fd_sc_hd__conb_1
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877__552 vssd1 vssd1 vccd1 vccd1 _10877__552/HI net552 sky130_fd_sc_hd__conb_1
X_08056_ net453 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ net390 _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a221o_1
X_05268_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ net423 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07007_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ _02649_ _02667_ _02668_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05199_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00912_ sky130_fd_sc_hd__xor2_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_101_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08958_ _01223_ _01413_ net411 vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__a21o_1
XANTENNA__07501__A_N net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ net257 _03370_ _03463_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08889_ _00708_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ net479 vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__o21a_1
XANTENNA__06587__Y _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net664 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XANTENNA__05932__B _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__A2 _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ net526 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08646__A1 _01475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ clknet_leaf_64_wb_clk_i _00603_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06657__B1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06409__B1 _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05379__B _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05947__X _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05395__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ clknet_leaf_79_wb_clk_i _00220_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10147_ clknet_leaf_16_wb_clk_i net722 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_89_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10078_ clknet_leaf_45_wb_clk_i _00136_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_85_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07118__C_N net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06673__B _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06240_ _01851_ _01869_ _01902_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__and3b_1
XANTENNA__07121__Y _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06392__C _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06171_ net197 net91 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05122_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__or2_1
Xhold304 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\]
+ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold315 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\] vssd1 vssd1
+ vccd1 vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold337 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\] vssd1 vssd1
+ vccd1 vccd1 net1006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09930_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\] _01786_
+ net153 net1007 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__o31a_1
XANTENNA__06281__D1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05053_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00763_ vssd1 vssd1
+ vccd1 vccd1 _00784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold359 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_down vssd1
+ vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09861_ _00762_ _04712_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__or3b_1
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06179__A2 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] _04160_
+ net942 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__o21ai_1
X_09792_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_107_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__mux2_1
X_05955_ net156 net147 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__nand2_2
XANTENNA__07128__A1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07128__B2 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout279_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04906_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] vssd1
+ vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _04053_ _04084_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_124_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05886_ _00715_ _01575_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07625_ net142 _03079_ _03182_ _03077_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07556_ _02235_ _03108_ _03109_ _01703_ _03112_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06507_ net100 _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__nor2_1
X_07487_ net179 _01744_ _02151_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__or3_1
XFILLER_0_107_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06438_ _02088_ _02110_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06369_ _02037_ _02041_ _02034_ _02035_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ _02672_ _03605_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__inv_2
XANTENNA__08143__X _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08039_ _03572_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net389 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05927__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10001_ clknet_leaf_32_wb_clk_i _00021_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ net568 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_54_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ net509 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__05026__A_N net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10765_ clknet_leaf_66_wb_clk_i _00586_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10696_ clknet_leaf_65_wb_clk_i _00527_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10973__613 vssd1 vssd1 vccd1 vccd1 _10973__613/HI net613 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05396__Y _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06014__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05369__B1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10733__RESET_B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05740_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] _00773_ vssd1
+ vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__or2_1
XANTENNA__05572__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05671_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ net416 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__or3b_1
XANTENNA__07530__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07410_ _02999_ _03000_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08390_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\] _03864_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07341_ _02945_ _02950_ _02952_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07272_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06223_ net200 _01829_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__nor2_4
XFILLER_0_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06154_ net91 _01834_ _01832_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__o21ai_1
Xhold101 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\] vssd1
+ vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__A1 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold123 _00327_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__dlygate4sd3_1
X_05105_ net480 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ _00821_ _00817_ net973 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a32o_1
Xhold134 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck vssd1 vssd1
+ vccd1 vccd1 net803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06085_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] vssd1 vssd1 vccd1 vccd1
+ _01770_ sky130_fd_sc_hd__or3b_1
Xhold145 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\] vssd1 vssd1
+ vccd1 vccd1 net814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold156 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\] vssd1 vssd1
+ vccd1 vccd1 net836 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _01781_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
X_05036_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\]
+ _00767_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__nor3_1
Xhold178 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] vssd1 vssd1
+ vccd1 vccd1 net858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09844_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\] _04848_ net264
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07962__B _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09775_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__or4bb_1
XANTENNA__07681__C _03144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] _02650_
+ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06572__A2 _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06578__B net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07026__Y _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ net865 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__mux2_1
XANTENNA__05482__B _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__A1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05938_ _00754_ _01631_ net100 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_1_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _00707_ _04050_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05869_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] net176
+ _01547_ net156 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07608_ _01811_ net163 _01672_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06594__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08588_ net816 net735 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07042__X _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07539_ _02080_ _02129_ _02150_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a21o_2
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10550_ clknet_leaf_12_wb_clk_i _00418_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _04420_ _04422_ _04421_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10481_ clknet_leaf_28_wb_clk_i _00349_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06260__A1 _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout97_X net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07760__B2 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__X _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10817_ net492 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08068__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10748_ clknet_leaf_64_wb_clk_i _00578_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08473__C1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06009__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05826__A1 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ clknet_leaf_26_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[11\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10823__498 vssd1 vssd1 vccd1 vccd1 _10823__498/HI net498 sky130_fd_sc_hd__conb_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06787__C1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06910_ _02579_ _02580_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07890_ _03442_ _03443_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__nand2_1
XANTENNA__06003__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06841_ net211 _02511_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__nor2_1
XANTENNA__06031__X _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ net785 net241 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
X_06772_ net93 _02414_ _02416_ net109 _02443_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a221o_1
X_08511_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__inv_2
X_05723_ net1017 _00824_ _00825_ net1038 _01430_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a221o_1
X_09491_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04613_ _04616_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__nand3_1
XFILLER_0_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08442_ net457 _03915_ _03695_ _03694_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__o211a_1
X_05654_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] _01301_
+ _01362_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08373_ team_07_WB.instance_to_wrap.team_07.buttonPixel _03700_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__o21a_1
X_05585_ _01286_ _01289_ _01291_ _01281_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout144_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07324_ _02939_ _00973_ _01109_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10437__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07255_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout409_A _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06206_ _01851_ _01869_ _01876_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07186_ _02835_ _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10814__D team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06137_ net286 net131 net127 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06068_ _01750_ _01751_ _01753_ _01754_ _01752_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a221o_1
Xfanout400 net402 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
Xfanout411 _00017_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout422 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_4
XFILLER_0_10_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05019_ net275 net272 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__nor2_2
Xfanout433 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] vssd1 vssd1
+ vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06589__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_2
XANTENNA__07037__X _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] vssd1
+ vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_2
X_09827_ _00657_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nor2_1
Xfanout477 net478 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_2
Xfanout488 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06545__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ _04767_ _04786_ _04787_ net244 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a32o_1
X_08709_ _04126_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ _04115_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__mux2_1
X_09689_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ _04736_ _00655_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a31o_1
XANTENNA__05940__B net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07213__A _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08028__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ clknet_leaf_35_wb_clk_i net875 net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout84 _02177_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_4
Xfanout95 net97 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10533_ clknet_leaf_31_wb_clk_i _00401_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05939__Y _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06481__A1 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ clknet_leaf_27_wb_clk_i net742 net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_up
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10395_ clknet_leaf_17_wb_clk_i _00039_ net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07981__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11016_ net387 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10325__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08446__C1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05370_ net433 _00668_ _01067_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__o21a_2
Xclkbuf_leaf_35_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08461__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload10 clknet_leaf_81_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinv_4
Xclkload21 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__06472__A1 _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07040_ _02214_ _02258_ _02692_ _02694_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a22o_1
Xclkload32 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__inv_6
XANTENNA__07496__C _03055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload43 clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_70_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload54 clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload54/X sky130_fd_sc_hd__clkbuf_8
Xclkload65 clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__inv_16
Xclkload76 clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_73_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07793__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__and4_1
XFILLER_0_103_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07942_ _01068_ net158 _01653_ _01083_ _01699_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07873_ _01051_ net118 _03427_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__o21a_1
X_09612_ _04664_ _04684_ net1092 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__o21ai_1
X_06824_ net427 net144 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09543_ net895 net222 _04605_ net902 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__a22o_1
X_06755_ _00671_ _00985_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout359_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__B1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05706_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__or2_1
X_09474_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ net266 net288 net219 vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a211o_1
X_06686_ _02338_ _02345_ _02346_ _02355_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08425_ _03638_ _03641_ net465 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__or3b_1
XFILLER_0_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05637_ net417 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01350_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08356_ _03828_ _03829_ _03831_ _03629_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__o211a_1
XANTENNA__06872__A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05568_ net415 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ _00677_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload4 clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_8
XANTENNA__08988__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07307_ _02930_ _02933_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[0\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] _03642_
+ _03639_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06591__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05499_ net418 _00692_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05266__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ net124 _01936_ _02861_ _02873_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__nor4_1
XANTENNA__07660__B1 _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07169_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] net298 net297 team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\]
+ _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10180_ clknet_leaf_22_wb_clk_i _00190_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout230 _02984_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_4
Xfanout252 _01489_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
Xfanout263 _00746_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_4
Xfanout274 _00651_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07715__A1 _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout285 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[1\] vssd1
+ vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_4
Xfanout296 _00969_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_4
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05951__A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09142__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07494__A3 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10516_ clknet_leaf_12_wb_clk_i _00384_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10447_ clknet_leaf_51_wb_clk_i _00331_ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06006__B net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10378_ clknet_leaf_4_wb_clk_i _00037_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07954__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__B team_07_WB.instance_to_wrap.team_07.labelPixel\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06022__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__A1 _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06390__B1 _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06676__B _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06540_ _00747_ net271 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06471_ _02064_ _02144_ _02137_ _02142_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_138_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08210_ _03688_ _03685_ _03687_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__and3b_1
X_05422_ _01007_ _01134_ _01107_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__or3b_1
X_09190_ net206 _04406_ _04408_ net402 net941 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07140__X _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ net54 net52 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05353_ _00966_ _01048_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08072_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ _03576_ net454 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05284_ net424 net425 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07023_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] _00829_ net297 team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08974_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] net824
+ net445 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07925_ _03320_ _03476_ _03478_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a211o_1
Xhold27 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05474__C _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold38 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ _01678_ _03321_ _03326_ _01689_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06807_ _02468_ _02469_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07787_ _01056_ _01597_ _01604_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04999_ net39 net38 net10 net9 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__or4_1
X_09526_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ net267 _04641_ net289 net220 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a221o_1
X_06738_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ net425 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ net413 _01416_ _04589_ net287 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o31a_1
X_06669_ _02340_ _02341_ _02339_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09870__A1 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ _03808_ _03882_ net484 vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09388_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08339_ net472 _03639_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10301_ clknet_leaf_24_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[14\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10232_ clknet_leaf_71_wb_clk_i net450 net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ clknet_leaf_22_wb_clk_i _00173_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input37_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[3\]
+ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05384__C _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05952__Y _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05681__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06496__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ net386 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05399__Y _01112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10758__RESET_B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07120__B _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__B1 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06017__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10184__D net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10340__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07927__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__Y _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06023__Y team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05938__B1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05971_ net173 net154 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__nor2_4
XFILLER_0_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07710_ _01729_ _02277_ _03206_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__a211o_1
X_04922_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
X_08690_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01757_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__nand2_1
XANTENNA__07155__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07641_ _01722_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__nand2_1
XANTENNA__06902__A2 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07572_ net137 net105 net165 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_105_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09311_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06523_ net98 net93 _02176_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__or3b_1
X_09242_ net228 _04446_ _04447_ net407 net1132 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06454_ net263 _02030_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__nor2_2
XANTENNA__06666__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04935__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05405_ _00669_ _01020_ _01061_ _01069_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__o22a_1
X_09173_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04391_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and3_1
X_06385_ net128 _01676_ net164 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06418__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08124_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or2_1
XANTENNA__07030__B _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05336_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] _00669_ vssd1
+ vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08055_ net453 net449 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__and3b_1
XANTENNA__07965__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05267_ net421 _00671_ _00979_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07006_ _02651_ _02659_ _02664_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05198_ _00909_ _00910_ _00908_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07918__A1 _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10010__RESET_B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05916__D net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _04246_ net420 _04245_ vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
X_07908_ _03369_ _03462_ _03368_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__a21oi_1
X_08888_ _00708_ _01429_ _04209_ net1070 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__a22o_1
XANTENNA__06597__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07839_ _03393_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__inv_2
XANTENNA__06354__B1 _02027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ net525 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09509_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ _04591_ net289 net221 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10774__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ clknet_leaf_64_wb_clk_i _00602_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07221__A _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06409__A1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06409__B2 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10215_ clknet_leaf_82_wb_clk_i _00219_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07891__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ clknet_leaf_16_wb_clk_i net769 net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ clknet_leaf_46_wb_clk_i net790 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06300__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06345__B1 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__X team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10979_ net619 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06648__A1 _02080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__B2 _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07131__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06170_ _01839_ _01842_ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and3b_1
XFILLER_0_26_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05121_ _00833_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
Xhold305 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\] vssd1 vssd1
+ vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold316 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\] vssd1 vssd1
+ vccd1 vccd1 net1007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__dlygate4sd3_1
X_05052_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00655_ _00761_
+ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__and3_1
XANTENNA__06820__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06820__B2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09860_ _00652_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _00772_
+ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__or3_1
XFILLER_0_110_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08811_ _04161_ _04162_ net192 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__a21oi_1
X_09791_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] _04808_ _04811_
+ _04813_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__a22o_1
X_08742_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ net239 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05954_ net160 _01566_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08673_ _04080_ _04098_ _04084_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_124_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05885_ _01574_ _01575_ _00715_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a21o_1
XANTENNA__06210__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07624_ _01666_ _01734_ _02278_ _03120_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__o2bb2a_1
X_07555_ _01666_ _03077_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06506_ net277 net89 net88 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__and3_2
XFILLER_0_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07486_ _01715_ _02045_ _03046_ _01714_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__and4b_1
XFILLER_0_9_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04430_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__and3_1
X_06437_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06368_ net168 _02040_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__nand2_1
XANTENNA__06880__A _01615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09053__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08107_ net914 _02671_ net1099 vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a21oi_1
X_05319_ _01029_ _01020_ _01024_ _01031_ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__and4b_1
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09087_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04328_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06299_ _01401_ net437 net434 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08038_ net409 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net392 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a221o_1
XANTENNA__06811__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10000_ clknet_leaf_32_wb_clk_i _00020_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout87_A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ clknet_leaf_32_wb_clk_i _00029_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10931__580 vssd1 vssd1 vccd1 vccd1 _10931__580/HI net580 sky130_fd_sc_hd__conb_1
XFILLER_0_118_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10902_ net567 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XANTENNA__08746__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07503__X team_07_WB.instance_to_wrap.team_07.memGen.stageDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ net508 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10764_ clknet_leaf_60_wb_clk_i _00585_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10695_ clknet_leaf_65_wb_clk_i _00526_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07886__A _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08481__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06014__B net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06566__B1 _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ clknet_leaf_43_wb_clk_i net813 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06581__A3 _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06030__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05670_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ net416 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_102_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07530__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10828__503 vssd1 vssd1 vccd1 vccd1 _10828__503/HI net503 sky130_fd_sc_hd__conb_1
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07340_ _01175_ _02417_ _02951_ _00965_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07271_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a21oi_1
X_09010_ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06222_ net154 _01736_ _01828_ net200 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a31o_2
XANTENNA__07796__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07046__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06153_ net103 _01828_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold102 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08404__B _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold113 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__dlygate4sd3_1
X_05104_ net1024 _00824_ _00825_ net1022 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a22o_1
Xhold124 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _00106_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlygate4sd3_1
X_06084_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__nand2_1
Xhold146 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\] vssd1 vssd1
+ vccd1 vccd1 net837 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] _01780_
+ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__nand2_1
X_05035_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__or4bb_1
Xhold179 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__dlygate4sd3_1
X_09843_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ _04844_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__and3_1
XANTENNA__06557__B1 _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_A _03033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06986_ _00713_ _02648_ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__nor2_1
X_09774_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06572__A3 _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06578__C net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05937_ net94 net86 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__nand2_2
X_08725_ _04134_ _04137_ _04136_ vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08849__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08656_ _01249_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__and2_1
X_05868_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _01546_
+ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__and3_1
XANTENNA__06875__A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ net184 _02073_ _02744_ _02863_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a211oi_2
XANTENNA__05532__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08587_ net735 net140 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05799_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ _01486_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__nand3_1
XFILLER_0_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _03091_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07469_ _00706_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ net392 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _04418_ _04419_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10480_ clknet_leaf_28_wb_clk_i _00348_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09139_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04370_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06115__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05954__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07760__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10816_ clknet_leaf_0_wb_clk_i _00036_ _00066_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10747_ clknet_leaf_64_wb_clk_i _00577_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06009__B net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05826__A2 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10678_ clknet_leaf_33_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[10\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_113_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06025__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__Y _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ net429 _00694_ _02510_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__o21a_1
XANTENNA__07200__B2 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06771_ net109 _02416_ _02441_ net116 _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ _03966_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__nand2_2
X_05722_ net475 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09490_ net986 net204 _04620_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__o21a_1
X_08441_ net458 _03914_ _03676_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05653_ _01349_ _01364_ _01365_ _01347_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__a31o_1
XANTENNA__05514__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03847_ _00727_
+ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05584_ _01295_ _01296_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07323_ net423 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout137_A _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07254_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ _02896_ _02899_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07019__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06205_ _01878_ _01885_ net97 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07185_ _01732_ _02836_ _01725_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_121_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout304_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06136_ _01808_ _01810_ _01815_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__and4_1
XFILLER_0_83_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06778__B1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06067_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__nand2_1
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_2
XANTENNA__05450__B1 _01103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05018_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net285
+ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__nand2_2
Xfanout412 team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1 vccd1
+ net412 sky130_fd_sc_hd__buf_2
XFILLER_0_100_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout423 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06222__X _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout445 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06589__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 net456 sky130_fd_sc_hd__buf_2
X_09826_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\] _04833_ vssd1 vssd1
+ vccd1 vccd1 _04838_ sky130_fd_sc_hd__and4_1
Xfanout467 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] vssd1
+ vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_2
Xfanout478 net483 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_2
Xfanout489 net491 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_2
XANTENNA__10365__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] _04783_ vssd1
+ vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__or2_1
X_06969_ _02562_ _02631_ _02636_ _02639_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_5_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08708_ net259 _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] _04738_ _04739_
+ _04734_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__o211a_1
X_08639_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05014__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10601_ clknet_leaf_35_wb_clk_i _00465_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout85 _02177_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10532_ clknet_leaf_30_wb_clk_i _00400_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05949__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout96 _01601_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463_ clknet_leaf_13_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_select
+ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06481__A2 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05020__Y _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05387__C _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05955__Y _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ net640 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__05509__A_N net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload11 clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_67_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload22 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_6
XFILLER_0_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload33 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload33/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_75_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xclkload44 clknet_leaf_71_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__clkinv_4
Xclkload55 clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload66 clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_114_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload77 clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08990_ _04258_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07972__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07941_ net257 _03310_ _03324_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__nor3_1
XANTENNA__10388__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07872_ net284 _01115_ _03390_ _03394_ _03288_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a311o_1
XFILLER_0_103_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05881__X _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _04666_ _04683_ _04684_ _04664_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a32o_1
X_06823_ net95 _02471_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09542_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ net221 _04605_ net853 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__a22o_1
X_06754_ net214 _02418_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05705_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__nor2_1
XANTENNA__07488__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09473_ net945 net203 _04609_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__o21a_1
X_06685_ _02079_ net84 _02329_ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08424_ net473 _03640_ net467 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a21oi_2
X_05636_ _01348_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08355_ net471 _03631_ _03659_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05567_ _01278_ _01279_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07306_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a21oi_1
Xclkload5 clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_117_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ _03763_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05498_ net418 _00692_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07237_ _01743_ _02758_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07660__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07168_ net447 team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\] net394 vssd1
+ vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__and3_1
X_06119_ _01723_ _01797_ _01799_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07099_ _02739_ _02751_ _02752_ _02748_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout220 _04582_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout231 net233 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
Xfanout242 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_4
Xfanout253 net255 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_4
Xfanout264 _04805_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
XANTENNA__07176__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_4
Xfanout286 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[1\] vssd1
+ vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
Xfanout297 _00942_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
X_09809_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\] net264 _04826_
+ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__o21ba_1
XANTENNA__05951__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05015__Y _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07511__X _03070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10515_ clknet_leaf_29_wb_clk_i _00383_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07651__A1 _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10446_ clknet_leaf_50_wb_clk_i _00330_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10377_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07954__A2 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06611__C1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06303__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08221__C _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__B _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__B1 _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06470_ net281 _01621_ _02104_ _02100_ net260 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06142__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05421_ _01061_ _01079_ _01097_ _01103_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_138_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__B1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08140_ _02670_ net145 vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_1
X_05352_ _00669_ _00967_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ _03575_ net454 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__mux2_1
XANTENNA__07642__A1 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05283_ _00993_ _00995_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__nand2_1
X_07022_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] net299 _02676_ vssd1
+ vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_112_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09395__A1 _01425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08973_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] net801
+ net445 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
Xhold17 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__B _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07924_ _03313_ _03315_ net252 vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__o21ai_1
Xhold28 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10287__RESET_B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold39 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07855_ net269 _03294_ _03299_ _03300_ _03285_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__o32a_1
XANTENNA__06905__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06806_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _02467_ _02476_
+ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a21bo_1
X_04998_ net19 net8 net33 net30 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__or4_2
X_07786_ _01597_ _01604_ _01056_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07044__A _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _01420_ _04640_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__or3b_1
X_06737_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ net425 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09456_ net929 net202 _04600_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06668_ net99 _01616_ _02312_ _02332_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06133__A1 _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06883__A _01615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _03707_ _03709_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21ai_1
X_05619_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ net443 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
X_06599_ net253 _01720_ _02271_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _01475_ net230 _04548_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08338_ net469 net467 vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07633__A1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ _03739_ _03747_ _03723_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ clknet_leaf_24_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[13\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05011__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10231_ clknet_leaf_81_wb_clk_i net451 net301 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10162_ clknet_leaf_18_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[9\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10093_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[2\]
+ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08749__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05962__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07164__A3 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10995_ net635 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_57_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__X _03814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__A0 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07872__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10861__536 vssd1 vssd1 vccd1 vccd1 _10861__536/HI net536 sky130_fd_sc_hd__conb_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07624__B2 _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold509 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10429_ clknet_leaf_21_wb_clk_i _00313_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07927__A2 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05938__A1 _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06033__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05970_ net256 _01657_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04921_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07640_ _01645_ _02744_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07571_ _01680_ net165 _01739_ _01685_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09310_ net225 _04493_ _04495_ net401 net1083 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06522_ net96 net89 _02176_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__nand2_1
X_06453_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] _02030_
+ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07863__B2 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05404_ _01057_ _01059_ _01070_ _00967_ _01116_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04391_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06384_ _01675_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_127_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\]
+ _03609_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__or2_1
XANTENNA__06418__A2 _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05335_ _00668_ net431 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__nor2_4
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07030__C _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ net1129 net293 _03580_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__a21o_1
X_05266_ net424 net425 _00978_ _00975_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ _02660_ _02664_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10468__RESET_B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05197_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00910_ sky130_fd_sc_hd__nand2_1
XANTENNA__07918__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ net474 net420 vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07907_ _01057_ net172 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__nand2_1
X_08887_ _03591_ _03592_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__mux2_2
XANTENNA__06597__B _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07838_ net272 _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__or2_1
XANTENNA__06354__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _03316_ _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ net220 _04605_ net868 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a22o_1
XANTENNA__05006__B net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10780_ clknet_leaf_64_wb_clk_i _00601_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09439_ net217 _04587_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06118__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05022__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05957__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07082__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06405__X _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10214_ clknet_leaf_79_wb_clk_i _00218_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10145_ clknet_leaf_15_wb_clk_i net758 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10076_ clknet_leaf_61_wb_clk_i _00134_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06345__A1 _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09295__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978_ net618 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_58_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07131__B net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06028__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05120_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold306 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold317 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold328 team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\] vssd1 vssd1 vccd1
+ vccd1 net997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold339 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\] vssd1 vssd1
+ vccd1 vccd1 net1008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05051_ _00781_ _00782_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\]
+ _00766_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[6\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08810_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] _04160_
+ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09790_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] _04810_ vssd1
+ vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08741_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__mux2_1
X_05953_ net178 _01645_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_107_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05884_ _01574_ _01575_ _00715_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a21oi_1
X_08672_ _04092_ _04089_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_124_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07623_ _02067_ _02150_ _03149_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10948__588 vssd1 vssd1 vccd1 vccd1 _10948__588/HI net588 sky130_fd_sc_hd__conb_1
X_07554_ net141 _03077_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06505_ _02109_ _02163_ _02169_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07485_ _01903_ _02040_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09224_ net228 _04433_ _04434_ net406 net1144 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09038__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06436_ _01680_ net167 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__and2_2
XFILLER_0_134_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09155_ net206 _04382_ _04383_ net401 net1113 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__a32o_1
X_06367_ net132 net122 net168 net142 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08106_ net914 _02671_ vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05318_ net190 _01014_ _01021_ _01030_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__o31a_1
XANTENNA__05777__A _01475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06298_ net177 _01973_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09086_ net208 _04331_ _04332_ net397 net1066 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06272__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08037_ net453 net449 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and3b_1
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05249_ _00957_ _00958_ _00961_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09988_ clknet_leaf_31_wb_clk_i _00027_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_08939_ net489 _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10901_ net566 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_84_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10832_ net507 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07232__A _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10763_ clknet_leaf_60_wb_clk_i _00584_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ clknet_leaf_69_wb_clk_i _00525_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05958__Y _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06566__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ clknet_leaf_43_wb_clk_i _00166_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06311__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ clknet_leaf_61_wb_clk_i _00117_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06030__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910__654 vssd1 vssd1 vccd1 vccd1 net654 _10910__654/LO sky130_fd_sc_hd__conb_1
XFILLER_0_78_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_29_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_102_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10867__542 vssd1 vssd1 vccd1 vccd1 _10867__542/HI net542 sky130_fd_sc_hd__conb_1
XANTENNA__07530__A3 _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06029__Y _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07270_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06221_ net176 net156 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06152_ _01644_ net103 net194 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07046__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold103 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
X_05103_ net475 _00814_ _00822_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__and3_2
Xhold114 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06083_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__or2_1
Xhold125 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\] vssd1 vssd1
+ vccd1 vccd1 net794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\] vssd1 vssd1
+ vccd1 vccd1 net805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold147 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\]
+ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09911_ net872 net152 net150 _04894_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a22o_1
X_05034_ _00763_ _00765_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__nand2_2
Xhold169 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\] vssd1
+ vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09842_ net1105 _04847_ _04849_ _04824_ vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__o22a_1
XANTENNA__06557__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06221__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\] _01769_ _04797_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] vssd1 vssd1 vccd1 vccd1
+ _04798_ sky130_fd_sc_hd__or4b_1
XFILLER_0_77_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06985_ _02647_ _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08724_ _01240_ _04080_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__and2_1
X_05936_ net115 net108 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__nand2_2
XANTENNA__06309__A1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _04073_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout451_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05867_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] net159
+ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07606_ _03078_ _03164_ _03159_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08586_ net145 _04027_ _03965_ vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__a21o_1
X_05798_ _01490_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_76_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07537_ net123 net143 _03079_ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__or4b_1
XANTENNA__07809__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__B2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ net291 _03035_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[29\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09207_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_119_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06493__B1 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06419_ _02074_ _02092_ _02090_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a21o_1
XANTENNA__07690__C1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05003__C net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ _02992_ _02993_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09138_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04369_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o31a_1
XFILLER_0_122_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09069_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ _04318_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05794__X _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05954__B _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06131__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05970__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input12_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06720__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10815_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.recHEART.heartDetect
+ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.heartPixel sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10746_ clknet_leaf_63_wb_clk_i _00576_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10096__Q team_07_WB.instance_to_wrap.team_07.labelPixel\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10677_ clknet_leaf_33_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[9\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07863__A1_N net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06025__B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A2 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06041__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _02417_ _02440_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__nand2_1
XANTENNA__06976__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05880__A _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05721_ net480 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ _00822_ _00824_ net973 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ _00731_ _03913_ _03679_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a21oi_1
X_05652_ _01331_ _01337_ _01342_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__or3b_1
XANTENNA__06711__A1 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08371_ _03777_ _03779_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__a21oi_1
X_05583_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] vssd1 vssd1 vccd1
+ vccd1 _01296_ sky130_fd_sc_hd__or3b_2
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07322_ _00672_ _02938_ _02937_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[0\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07267__A2 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07253_ _00718_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06204_ net94 _01879_ _01883_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07184_ _01715_ _01873_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__nor2_4
XFILLER_0_108_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_wb_clk_i_X clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06135_ net280 _01812_ _01813_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06066_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05017_ _00635_ _00649_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__nor2_1
Xfanout402 net405 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
Xfanout413 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_4
Xfanout435 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[2\] vssd1 vssd1 vccd1
+ vccd1 net435 sky130_fd_sc_hd__buf_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_2
XANTENNA_input4_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ net1075 _04834_ _04837_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__o21a_1
XANTENNA__07047__A _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] vssd1 vssd1
+ vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_2
Xfanout468 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[2\] vssd1
+ vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_2
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_2
X_09756_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] _04783_ vssd1
+ vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__nand2_1
XANTENNA__06886__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ _02556_ _02637_ _02638_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a21o_1
X_08707_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ _01238_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__a41o_1
X_05919_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] _01593_
+ _01580_ _01578_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__o2bb2a_1
X_09687_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] _04738_ vssd1
+ vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06899_ net286 _02568_ _02562_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_90_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10963__603 vssd1 vssd1 vccd1 vccd1 _10963__603/HI net603 sky130_fd_sc_hd__conb_1
X_08638_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ net455 _04062_ _04063_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__o311a_1
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08569_ _04015_ _04016_ _03996_ vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10600_ clknet_leaf_34_wb_clk_i _00464_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05014__B net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout86 _01629_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10531_ clknet_leaf_31_wb_clk_i _00399_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout97 _01601_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ clknet_leaf_27_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_up
+ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10393_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[1\]
+ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05965__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06413__X _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11014_ net386 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05971__Y _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_X net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10729_ clknet_leaf_59_wb_clk_i _00559_ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload12 clknet_leaf_83_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_8
Xclkload23 clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_6
XANTENNA__06036__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload34 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__bufinv_16
Xclkload45 clknet_leaf_72_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload45/X sky130_fd_sc_hd__clkbuf_4
Xclkload56 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_114_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload67 clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_16
Xclkload78 clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_114_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05875__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ _01067_ net216 _03314_ _03494_ net252 vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_110_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06042__Y _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10916__660 vssd1 vssd1 vccd1 vccd1 net660 _10916__660/LO sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_44_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07871_ _03421_ _03422_ _03340_ _03346_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__a211o_1
XANTENNA__07185__A1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] _04682_ vssd1
+ vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__nand2_1
X_06822_ net95 _02471_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__and2_1
X_09541_ _04651_ net853 net220 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
X_06753_ _00973_ net198 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__nor2_1
X_05704_ net413 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01415_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__or3_1
X_09472_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ net266 net288 net219 vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a211o_1
XANTENNA__07488__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06684_ _02336_ _02349_ _02352_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__and3b_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08423_ net768 _03897_ net129 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05635_ net416 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01348_ sky130_fd_sc_hd__and3b_1
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08354_ _03632_ _03637_ _03766_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08437__A1 _00711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05566_ _01270_ _01272_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__xnor2_1
X_07305_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_22_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ net466 _03641_ _03660_ _03667_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__o311a_1
X_05497_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01201_ _01208_ _01209_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__or4b_1
Xclkload6 clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07236_ net169 _02082_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07660__A2 _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] net299 _02673_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06118_ net197 _01798_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__nand2_1
X_07098_ net143 _01669_ _01664_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a21o_1
X_06049_ net176 _01737_ net179 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__o21ai_1
Xfanout210 net213 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_4
Xfanout221 _04582_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
Xfanout243 _04824_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_1
Xfanout265 _04591_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
XANTENNA__07176__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 _00650_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
Xfanout287 _04584_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_4
X_09808_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\] _04825_ vssd1
+ vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__and2_1
Xfanout298 _00831_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06923__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09739_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] _04772_ vssd1
+ vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05025__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10514_ clknet_leaf_12_wb_clk_i _00382_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08770__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07651__A2 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05966__Y _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ clknet_leaf_41_wb_clk_i _00329_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__B1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[1\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06611__B1 _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05982__X _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10401__SET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__A2 _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09987__D net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05420_ _01026_ _01110_ _01132_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07150__A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05351_ net431 net393 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__nor2_2
XFILLER_0_138_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08070_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ net392 _03026_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ _03588_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__a221o_1
X_05282_ _00994_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07021_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] net298 net297 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\]
+ _02675_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05876__Y _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06401__A_N _02074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] net840
+ net445 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
X_07923_ _03312_ _03477_ _03317_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__a21oi_1
Xhold18 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__C net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold29 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ _03364_ _03389_ _03402_ _03403_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06805_ _02466_ _02467_ _02468_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__or3_1
X_07785_ _01115_ net110 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04997_ net35 net34 net37 net36 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__or4_1
X_09524_ _00665_ _00666_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__nor2_1
X_06736_ _02406_ _02407_ _02408_ _02326_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recHEART.heartDetect
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09455_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ net265 _04599_ net287 net217 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
X_06667_ _02108_ _02312_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__nor2_1
X_08406_ _03709_ _03880_ _03742_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__o21a_1
X_05618_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] _01327_
+ _01330_ _01324_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__o211a_1
X_09386_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _01424_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__nor2_1
X_06598_ net251 _02270_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__nor2_2
X_08337_ _03715_ _03813_ _03752_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_35_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05549_ _01259_ _01261_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08268_ _03709_ _03746_ _03742_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _02856_ _02860_ _01744_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a21oi_1
X_08199_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\] _01255_ vssd1
+ vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ clknet_leaf_75_wb_clk_i _00041_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10161_ clknet_leaf_18_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[8\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10092_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[1\]
+ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07506__Y _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05962__B _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08765__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ net634 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10378__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07085__B1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10902__567 vssd1 vssd1 vccd1 vccd1 _10902__567/HI net567 sky130_fd_sc_hd__conb_1
XFILLER_0_122_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10428_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[2\]
+ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06045__D1 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10359_ clknet_leaf_3_wb_clk_i net714 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06033__B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06060__A1 _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04920_ net3 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_109_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07145__A _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06036__D_N _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ _02208_ _03126_ _03127_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06521_ _02088_ _02194_ _01646_ _01739_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__or2_1
X_06452_ _02125_ _02123_ _02122_ _02121_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__and4b_1
XFILLER_0_29_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05403_ net190 _01025_ _01102_ _01068_ _01038_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__o32a_1
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ net207 _04393_ _04394_ net403 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06383_ _01675_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__or2_1
X_05334_ net421 _01046_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__and2_1
XANTENNA__06418__A3 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08053_ net448 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net389 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05265_ _00975_ _00977_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout112_A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07004_ _00713_ _02666_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05196_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00909_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06224__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08955_ net474 _00827_ _01431_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_129_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout481_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ _03373_ _03459_ _03460_ _03457_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08879__A1 _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ net435 _04208_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__xnor2_1
X_07837_ _03288_ _03351_ _03390_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__nand3b_1
XANTENNA__07551__A1 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10090__RESET_B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _01083_ net183 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09507_ net868 net204 _04631_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06719_ _02390_ _02391_ _02389_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a21bo_1
X_10884__559 vssd1 vssd1 vccd1 vccd1 _10884__559/HI net559 sky130_fd_sc_hd__conb_1
XFILLER_0_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ net108 _03253_ _03254_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09438_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01415_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ net224 _04535_ _04536_ net397 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05022__B _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05957__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10213_ clknet_leaf_72_wb_clk_i _00217_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_37_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input42_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05973__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ clknet_leaf_15_wb_clk_i net723 net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_10819__494 vssd1 vssd1 vccd1 vccd1 _10819__494/HI net494 sky130_fd_sc_hd__conb_1
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10075_ clknet_leaf_61_wb_clk_i _00133_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07542__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06345__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06750__C1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10977_ net617 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__10232__SET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05867__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] vssd1 vssd1
+ vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_back vssd1
+ vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
X_05050_ _00776_ _00775_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold329 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] vssd1 vssd1
+ vccd1 vccd1 net998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05883__A _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ net1117 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__mux2_1
X_05952_ net178 _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_4
XANTENNA__06050__Y _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08671_ _04096_ _04097_ net1165 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__a21o_1
X_05883_ _01574_ _01575_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_124_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07622_ _03119_ _03179_ _03176_ _03170_ _03168_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_124_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07553_ _01660_ _03080_ _03111_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a21oi_1
X_06504_ _02148_ _02176_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__nand2_2
X_07484_ _02278_ _03042_ _03043_ _01659_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04430_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05123__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06435_ net273 _00753_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__and2_4
XFILLER_0_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07049__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__or2_1
XANTENNA__10017__SET_B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06366_ _01651_ _01698_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__nor2_4
XANTENNA__06506__X _02180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08105_ net803 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs _00244_
+ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05317_ net188 _01004_ _01014_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09085_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04328_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout115_X net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06297_ net434 _01396_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__or2_1
XANTENNA__06225__Y _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ _03570_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net389 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05248_ net491 _00797_ _00960_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05179_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00886_ vssd1 vssd1
+ vccd1 vccd1 _00892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09987_ clknet_leaf_33_wb_clk_i net411 net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07772__B2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\] _04234_
+ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__and2_1
XANTENNA__07509__D1 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ net258 _04192_ _04197_ _04195_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__a31o_1
XFILLER_0_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10900_ net565 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_4_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10831_ net506 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10762_ clknet_leaf_66_wb_clk_i _00583_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10693_ clknet_leaf_69_wb_clk_i _00524_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05968__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06263__A1 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07212__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10127_ clknet_leaf_43_wb_clk_i _00165_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07407__B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10058_ clknet_leaf_61_wb_clk_i net807 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07515__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06039__A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10908__573 vssd1 vssd1 vccd1 vccd1 _10908__573/HI net573 sky130_fd_sc_hd__conb_1
XFILLER_0_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06220_ _01868_ _01871_ _01854_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06151_ net95 _01831_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07046__A3 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05102_ net475 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ _00822_ _00824_ net968 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a32o_1
Xhold104 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
X_06082_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] _01766_ _01761_
+ _01748_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold126 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold137 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[6\] vssd1 vssd1
+ vccd1 vccd1 net806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09910_ _01780_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05033_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\]
+ _00764_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__o21ai_1
Xhold159 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09841_ _00657_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nor2_1
XANTENNA__06557__A2 _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] vssd1 vssd1 vccd1 vccd1
+ _04797_ sky130_fd_sc_hd__nand3_1
X_06984_ _00712_ _00714_ _02645_ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__or3b_1
XANTENNA__06221__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ _04034_ _04082_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__a31o_1
X_05935_ net118 net111 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout277_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ _04079_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__or2_1
X_05866_ _01552_ _01556_ _01553_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a21oi_2
XANTENNA__04957__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07605_ net155 net107 _03161_ _03163_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08585_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ _03622_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05797_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _01485_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] vssd1 vssd1
+ vccd1 vccd1 _01491_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout444_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07536_ _02223_ _03093_ _03094_ _01612_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07467_ net409 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net391 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09206_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06418_ net107 _01697_ net164 _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a31o_2
XFILLER_0_9_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06493__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07690__B1 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _02990_
+ net476 vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06349_ net414 net135 _02016_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__o31a_1
XFILLER_0_115_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08019_ net1138 net40 net42 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__and3b_1
XFILLER_0_124_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout92_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06131__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06181__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08058__B net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06720__A2 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10814_ clknet_leaf_58_wb_clk_i team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect
+ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.playButtonPixel
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08773__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10745_ clknet_leaf_62_wb_clk_i _00575_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10676_ clknet_leaf_33_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[8\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06236__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07984__A1 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06787__A2 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A3 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06041__B _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06976__B _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05720_ net1061 _00824_ _00825_ net969 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__a22o_1
XANTENNA__05880__B _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05651_ _01352_ _01354_ _01357_ _01363_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06711__A2 _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08370_ net487 _00727_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05582_ _01286_ _01292_ _01294_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07321_ net424 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ _02898_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07672__B1 _02081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06203_ net94 _01879_ _01880_ net109 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07183_ net159 _01699_ _01718_ _01829_ net201 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o311a_2
XFILLER_0_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06134_ _01812_ _01813_ net280 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06065_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05016_ net285 net284 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__nand2_1
Xfanout403 net405 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_2
XFILLER_0_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout414 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col vssd1 vssd1
+ vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07727__A1 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout425 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout394_A _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout436 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 net436 sky130_fd_sc_hd__clkbuf_2
Xfanout447 team_07_WB.instance_to_wrap.team_07.memGen.stage\[0\] vssd1 vssd1 vccd1
+ vccd1 net447 sky130_fd_sc_hd__buf_2
X_09824_ _04827_ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nor2_1
XANTENNA__07047__B net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\] vssd1 vssd1
+ vccd1 vccd1 net458 sky130_fd_sc_hd__buf_2
Xfanout469 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[2\] vssd1
+ vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09755_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] _04783_ vssd1
+ vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and2_1
X_06967_ net105 _02497_ _02543_ _02627_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout182_X net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__A2 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05918_ net100 net87 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__or2_1
X_08706_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ _04121_ _04124_ _04115_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__o22a_1
X_09686_ net1139 _04735_ _04737_ _04730_ _04734_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__o221a_1
X_06898_ net270 _02568_ _02562_ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08637_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__xnor2_1
X_05849_ _01538_ _01542_ _01536_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_7_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08568_ net54 net52 net139 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07519_ _01873_ _02744_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08499_ _03964_ _03965_ vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10530_ clknet_leaf_31_wb_clk_i _00398_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout87 _01610_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_4
XFILLER_0_107_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout98 net99 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06407__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10461_ clknet_leaf_29_wb_clk_i net1014 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10392_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[2\]
+ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07966__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07238__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07718__A1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ net387 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08768__S net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05901__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10728_ clknet_leaf_59_wb_clk_i _00558_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10659_ clknet_leaf_19_wb_clk_i _00514_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload13 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10374__RESET_B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload24 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_12
XFILLER_0_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload35 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__bufinv_16
Xclkload46 clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_8
Xclkload57 clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_114_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload68 clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__inv_16
Xclkload79 clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__inv_6
XANTENNA__05875__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09159__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06052__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__B1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _03361_ _03424_ _03419_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07185__A2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ net92 _02467_ _02474_ _02491_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__o31ai_1
X_10986__626 vssd1 vssd1 vccd1 vccd1 _10986__626/HI net626 sky130_fd_sc_hd__conb_1
X_09540_ _01419_ net289 _04645_ net267 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a32o_1
X_06752_ net424 _00981_ net183 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_13_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09331__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05703_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01415_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__nor2_1
X_09471_ net920 net202 _04608_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__o21a_1
XANTENNA__07456__A_N net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06683_ _02345_ _02346_ _02355_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__and3_1
X_08422_ _03894_ _03896_ _03888_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__o21a_1
X_05634_ net440 _01280_ _01327_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08353_ _03760_ _03825_ _03827_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a31o_1
X_05565_ _01274_ _01277_ _01276_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__or3b_2
XFILLER_0_117_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout142_A _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07304_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08284_ net472 _03761_ _03760_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_12
X_05496_ net418 _00690_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07235_ _02876_ _02879_ _02881_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__o31a_1
XFILLER_0_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07660__A3 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07166_ _02799_ _02816_ _02818_ _02806_ _02814_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\]
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04970__A team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07948__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06117_ net181 _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__nand2_2
XANTENNA__07948__B2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08070__B1 _03026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07097_ _02138_ net82 _02732_ _02750_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a22o_1
XANTENNA__05959__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06048_ net160 _01735_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nor2_2
Xfanout200 _01662_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_4
Xfanout211 net213 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
Xfanout222 _04582_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_2
Xfanout233 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout244 _04765_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
Xfanout255 _01488_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_2
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout266 _04591_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_2
X_09807_ net243 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__inv_2
Xfanout277 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
Xfanout288 _04584_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
Xfanout299 _00829_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06384__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__xor2_1
X_09738_ _04767_ _04771_ _04773_ net245 net1035 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09669_ _04716_ _04725_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_16_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07521__A _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06408__Y _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__RESET_B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ clknet_leaf_29_wb_clk_i _00381_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05976__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10444_ clknet_leaf_49_wb_clk_i _00328_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07939__A1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ clknet_leaf_2_wb_clk_i net691 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06611__A1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06611__B2 _02282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06375__B1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05717__A3 _01425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07415__B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07150__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05350_ _01062_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06047__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05281_ _00976_ _00978_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07020_ net394 _02674_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06334__X _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08971_ net415 net817 net445 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
X_07922_ _01067_ net172 vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__nand2_1
Xhold19 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _03379_ _03404_ _03406_ _03407_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06510__A _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ net92 _02474_ _02471_ net95 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__o2bb2a_1
X_07784_ _01058_ net108 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nand2_1
X_04996_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\] vssd1 vssd1
+ vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ net891 net205 _04639_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__o21a_1
X_06735_ _02311_ _02356_ _01413_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout357_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _04598_ _04597_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__o21ai_1
X_06666_ net98 _01616_ _02312_ net274 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08405_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03879_ _00727_
+ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__o21a_1
X_05617_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01319_
+ _01325_ _01315_ _01329_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__o221a_1
X_09385_ _00659_ _04546_ _04547_ _04542_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06597_ net157 _02021_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08336_ net462 _03803_ _03812_ _03797_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05548_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] vssd1 vssd1 vccd1
+ vccd1 _01261_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08871__S net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08291__B1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ net412 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03745_
+ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__nor3_1
XFILLER_0_62_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05479_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared _01191_ vssd1 vssd1
+ vccd1 vccd1 _01192_ sky130_fd_sc_hd__or2_2
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07633__A3 _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04971__Y _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ _01645_ _01734_ _02867_ _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06244__X _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08198_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\] _01379_ vssd1
+ vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__nand2_1
X_07149_ _02800_ _02801_ _02798_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__o21a_1
X_10160_ clknet_leaf_18_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10091_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[0\]
+ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09543__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08111__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10993_ net633 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_96_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07085__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10427_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[1\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06045__C1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10358_ clknet_leaf_1_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear
+ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.maze_clear_edge_detector.inter
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06060__A2 _01481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ clknet_leaf_42_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[2\]
+ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06330__A team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06520_ net201 _02089_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__or2_2
XANTENNA__05233__X _00946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06451_ net167 _01711_ _01734_ _02058_ _02092_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06048__Y _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05402_ net393 _01058_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__nand2_2
X_09170_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04391_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06382_ net178 _01873_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__or2_4
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08121_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05333_ _00966_ net296 _01045_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_126_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08052_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ net294 _03579_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05264_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _00973_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07003_ _02649_ _02665_ _02648_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05195_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00901_ vssd1 vssd1
+ vccd1 vccd1 _00908_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06224__B _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout105_A _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08954_ net490 _00797_ _01427_ _01428_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_129_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07905_ net257 _03382_ _03385_ _03386_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__nor4_1
X_08885_ _04205_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout474_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07055__B _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ _03390_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__inv_2
XANTENNA__07551__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04979_ net472 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
X_07767_ _01084_ net187 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09506_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ net268 net290 net220 vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06718_ _02066_ _02313_ net83 _02170_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22oi_1
X_07698_ net273 net93 net115 _01609_ _02009_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06649_ _02127_ _02297_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__nand2_1
X_09437_ net413 _01414_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10999__636 vssd1 vssd1 vccd1 vccd1 _10999__636/HI net636 sky130_fd_sc_hd__conb_1
X_09368_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04533_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07067__B2 _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ net411 net462 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nor2_1
X_09299_ net979 net396 net225 _04487_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06814__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10212_ clknet_leaf_72_wb_clk_i _00216_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05973__B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ clknet_leaf_15_wb_clk_i net715 net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_89_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input35_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ clknet_leaf_61_wb_clk_i _00132_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07542__A2 _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08077__A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ net616 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_63_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06325__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold308 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\] vssd1
+ vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold319 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] vssd1 vssd1
+ vccd1 vccd1 net988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06281__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06569__B1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07230__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05883__B _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05951_ net180 net176 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__nand2_4
X_08670_ _04054_ _04058_ _04073_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05882_ _01574_ _01575_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07621_ _03177_ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ _01739_ net163 _03110_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06503_ _02148_ _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07483_ _02278_ _03042_ _03043_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__o21ai_1
X_09222_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04430_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__nand2_1
X_06434_ net262 _02030_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__or2_4
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08715__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__nand2_1
XANTENNA__07049__A1 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06365_ _02034_ _02035_ _02038_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08104_ net762 net759 _02671_ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05316_ _01026_ _01028_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__or2_1
X_09084_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04328_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__nand2_1
X_06296_ net160 _01969_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08035_ net409 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net291 _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a221o_1
X_05247_ _00683_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared vssd1
+ vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout108_X net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05178_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00890_ vssd1 vssd1
+ vccd1 vccd1 _00891_ sky130_fd_sc_hd__xnor2_1
X_09986_ clknet_leaf_79_wb_clk_i _00091_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_10851__526 vssd1 vssd1 vccd1 vccd1 _10851__526/HI net526 sky130_fd_sc_hd__conb_1
XANTENNA__07066__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ _01432_ _01484_ _01762_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__and3_2
XANTENNA__07509__C1 _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ net297 _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07819_ _01057_ net171 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08799_ _04153_ _04154_ net192 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__a21oi_1
X_10830_ net505 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05314__A _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10761_ clknet_leaf_62_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\]
+ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ clknet_leaf_68_wb_clk_i _00523_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05968__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05984__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06432__X _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07212__A1 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10126_ clknet_leaf_43_wb_clk_i _00164_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10399__RESET_B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05990__Y _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05208__B _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ clknet_leaf_61_wb_clk_i _00115_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07515__A2 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07704__A _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload0_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05224__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10959_ net599 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_70_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05230__Y _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06150_ net181 net177 _01657_ net103 _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a41o_1
XANTENNA__06055__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05101_ net479 team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00810_ _00816_
+ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__and4_2
XFILLER_0_130_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06081_ _01762_ _01767_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__or2_1
Xhold105 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\] vssd1 vssd1
+ vccd1 vccd1 net774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold127 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _00116_ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
X_05032_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__nor2_1
Xhold149 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[2\]
+ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08270__A _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] _04844_ vssd1
+ vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06502__B net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954__594 vssd1 vssd1 vccd1 vccd1 _10954__594/HI net594 sky130_fd_sc_hd__conb_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ _04796_ _04794_ net1004 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06983_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] _02645_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] vssd1 vssd1
+ vccd1 vccd1 _02647_ sky130_fd_sc_hd__a21o_1
X_08722_ _04135_ _04134_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__mux2_1
X_05934_ net116 _01616_ _01626_ _01610_ _01600_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__a311oi_4
XTAP_TAPCELL_ROW_1_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05865_ _01547_ net156 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__nand2_1
X_08653_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01239_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or3_1
XANTENNA__06714__B1 _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07604_ net138 _01688_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05796_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] _01486_
+ _01487_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__and3_1
XANTENNA__06190__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08584_ net145 _04026_ _03965_ vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07535_ net100 _02107_ _02191_ _03072_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__o31a_1
XFILLER_0_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout437_A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net292 _03034_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[28\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA__06517__X _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09205_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06417_ net214 net173 _01698_ _01684_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06493__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08219__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _02990_
+ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07690__B2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06348_ _02012_ _02022_ _02019_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__or3b_1
X_09136_ net4 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ _04368_ vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
X_09067_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ net6 _04317_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
X_06279_ _01662_ _01954_ _01955_ _01952_ _01944_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08018_ net987 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_back
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10892__648 vssd1 vssd1 vccd1 vccd1 net648 _10892__648/LO sky130_fd_sc_hd__conb_1
XFILLER_0_124_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06548__A3 _02180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05309__A _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ clknet_leaf_72_wb_clk_i _00074_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06131__C _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07524__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10813_ clknet_leaf_59_wb_clk_i _00634_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10100__D team_07_WB.instance_to_wrap.team_07.memGen.stageDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10744_ clknet_leaf_63_wb_clk_i _00574_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07130__B1 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06427__X _02101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ clknet_leaf_33_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[7\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05985__Y _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07984__A2 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ clknet_leaf_52_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireHighlightDetect
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05650_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] _01301_
+ _01362_ _01360_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06172__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05581_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01253_
+ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07320_ _01190_ _01192_ _01193_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07251_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ _02897_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07672__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07672__B2 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06202_ net109 _01880_ _01881_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07182_ _02134_ net82 _02741_ _02831_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06133_ _01812_ _01813_ net280 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08712__B net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07609__A _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06064_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05015_ _00649_ net275 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__nor2_4
XFILLER_0_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
XANTENNA__07188__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout415 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] vssd1
+ vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_2
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07727__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout426 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09823_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] _04834_ vssd1
+ vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__and2_1
Xfanout437 net438 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout448 net450 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_2
XANTENNA__07047__C _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout459 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\] vssd1 vssd1
+ vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
X_09754_ net965 _04782_ _04784_ net244 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__o22a_1
X_06966_ _02488_ _02560_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__nand2_1
XANTENNA__07344__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ _04122_ _04123_ net242 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__a21oi_1
X_05917_ net89 net88 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__nand2_2
X_09685_ _04730_ _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06897_ _02549_ _02567_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08636_ _00693_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__or2_1
X_05848_ _01540_ _01541_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08567_ _03615_ _04014_ net139 vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a21oi_1
X_05779_ _01468_ _01471_ _01473_ _01459_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07518_ net179 _01657_ net256 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_65_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08498_ _02670_ net145 _03652_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nor3_2
XFILLER_0_130_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07449_ net451 net448 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__and2_2
Xfanout88 _01609_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_4
Xfanout99 _01600_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_4
XFILLER_0_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10460_ clknet_leaf_27_wb_clk_i net1028 net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09119_ net209 _04354_ _04356_ net400 net1021 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__a32o_1
X_10391_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[1\]
+ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07966__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857__532 vssd1 vssd1 vccd1 vccd1 _10857__532/HI net532 sky130_fd_sc_hd__conb_1
XFILLER_0_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08114__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07238__B _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] vssd1 vssd1 vccd1
+ vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout88_X net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__A2 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ net639 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XANTENNA__05981__B _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05326__X _01039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10388__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10727_ clknet_leaf_60_wb_clk_i _00557_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07654__A1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05221__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10658_ clknet_leaf_20_wb_clk_i _00513_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload14 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_24_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06036__C _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload25 clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_51_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload36 clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__08603__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload47 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinv_8
X_10589_ clknet_leaf_36_wb_clk_i _00453_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06604__Y _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload58 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__bufinv_16
Xclkload69 clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_114_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06052__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08959__S _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ net92 _02467_ _02477_ net113 _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__a221o_1
X_06751_ net424 _00981_ net183 _02420_ _02422_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a32o_1
XFILLER_0_92_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05702_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__or2_2
X_09470_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ net265 net287 net219 vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a211o_1
X_06682_ _02336_ _02339_ _02343_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__or3b_1
XFILLER_0_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07451__X _03026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08421_ _03656_ _03667_ _03895_ _03890_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__a31o_1
X_05633_ net439 _01322_ _01344_ _01345_ _01320_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_114_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08352_ _03760_ _03825_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_53_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_05564_ _01266_ _01270_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__nor2_1
XANTENNA__06508__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07303_ net441 _01328_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08283_ net466 _03643_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__nand2_1
X_05495_ net418 _00690_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06227__B _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinv_4
X_07234_ _02882_ _02884_ _02880_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07165_ net166 _02033_ _02758_ _02817_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06116_ net175 net123 _01702_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__or3_2
X_07096_ _01618_ _01921_ _02196_ net260 _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a221o_4
XANTENNA__05959__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06243__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06047_ net125 _01699_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__nand2_2
XFILLER_0_121_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10084__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 _01661_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_4
XFILLER_0_100_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_4
Xfanout223 _04510_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
XFILLER_0_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
Xfanout245 _04765_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_4
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
X_09806_ _04798_ _04804_ _04807_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09570__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06384__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_2
XFILLER_0_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07998_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__xor2_1
XANTENNA__07581__B1 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__inv_2
X_06949_ net174 _02506_ _02508_ _02581_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_69_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09668_ _04716_ _04724_ _04725_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__nor3_1
XANTENNA__07333__A0 _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08619_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__or2_1
X_09599_ _04665_ _04675_ net1142 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10928__577 vssd1 vssd1 vccd1 vccd1 _10928__577/HI net577 sky130_fd_sc_hd__conb_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07636__A1 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10512_ clknet_leaf_12_wb_clk_i _00380_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10443_ clknet_leaf_41_wb_clk_i net792 net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10374_ clknet_leaf_18_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[2\]
+ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06611__A2 _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05992__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__X _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06375__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05216__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09864__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07431__B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07627__A1 _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06047__B _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05280_ _00988_ _00992_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__nand2_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05886__B _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10524__RESET_B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08970_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] net821
+ net444 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
X_07921_ net132 net121 _03475_ _03473_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__a31o_1
X_07852_ net105 _03376_ _03387_ net106 vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06803_ net430 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1
+ vccd1 vccd1 _02474_ sky130_fd_sc_hd__xnor2_2
Xinput1 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
X_07783_ _03285_ _03286_ _03337_ _03336_ _03335_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__o32a_1
X_04995_ net458 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
X_09522_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ net267 _04638_ net220 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a211o_1
X_06734_ _02307_ _02359_ _01223_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09453_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] vssd1
+ vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__and2b_1
X_06665_ _02334_ _02336_ _02337_ _02330_ _02259_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout252_A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ _03745_ _03804_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__nor2_1
X_05616_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] net441
+ _01328_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__a21o_1
X_09384_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ net397 _04308_ net224 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06596_ _02267_ _02264_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08335_ _03718_ _03811_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__nor2_1
X_05547_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08266_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] _03744_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a21oi_1
X_05478_ _00795_ _00963_ net486 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07217_ net179 _02033_ _02863_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08197_ net458 _01381_ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__a21oi_1
X_07148_ _02072_ _02758_ _02781_ _02059_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07079_ _02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__inv_2
X_10090_ clknet_leaf_66_wb_clk_i _00148_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06701__A _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10992_ net632 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06148__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05987__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06435__X _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10426_ clknet_leaf_18_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[0\]
+ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06045__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10357_ clknet_leaf_56_wb_clk_i _00297_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10288_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[1\]
+ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07713__Y _03269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07848__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__B2 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06450_ net166 _01734_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08972__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06058__A _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05401_ _00970_ _01031_ _01089_ _01090_ _01101_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__o221a_1
X_06381_ net178 _01873_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05332_ _01018_ _01039_ _01044_ _01032_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__or4b_1
X_08120_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08273__A _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08051_ net449 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net390 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05263_ net424 net425 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__nand2_1
X_07002_ _02649_ _02664_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05194_ _00902_ _00903_ _00905_ _00906_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08953_ net491 _04243_ vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07904_ net154 _03374_ _03458_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__or3b_1
X_08884_ _01399_ _01397_ _04203_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07835_ net273 _01055_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ _03307_ _03319_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__nor2_1
X_04978_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs vssd1 vssd1 vccd1
+ vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs sky130_fd_sc_hd__inv_2
X_09505_ net908 net222 _04605_ net934 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ _02079_ _02258_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ net119 _02031_ _02148_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__and2b_1
X_06648_ _02080_ _02287_ _02289_ _02135_ _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__o221a_1
XFILLER_0_94_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09367_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04533_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__or2_1
X_06579_ _01627_ _02106_ _02149_ _02251_ _02252_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10446__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ _03722_ _03795_ _03718_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09298_ _04485_ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05078__B2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06814__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ net460 _01282_ _01308_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06415__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10211_ clknet_leaf_72_wb_clk_i _00215_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10142_ clknet_leaf_16_wb_clk_i _00042_ net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_37_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10073_ clknet_leaf_61_wb_clk_i _00131_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07527__B1 _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10103__D team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06750__A1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ net615 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10187__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06606__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold309 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] vssd1 vssd1
+ vccd1 vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10409_ clknet_leaf_1_wb_clk_i _00300_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07230__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06341__A _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05950_ net185 net171 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07518__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05881_ _01565_ _01573_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__or2_4
XFILLER_0_75_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08191__B1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _01721_ _03079_ _03120_ _01733_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_124_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07613__A2_N net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07551_ _01658_ net170 _01701_ _01669_ _01664_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__o32a_1
XFILLER_0_89_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06502_ _01582_ net115 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_17_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07482_ _01489_ net185 _01901_ _01664_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ net227 _04431_ _04432_ net406 net883 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06433_ net262 _02030_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__nor2_4
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08274__Y _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09152_ net206 _04380_ _04381_ net401 net933 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__a32o_1
X_06364_ net168 _02036_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08103_ net761 _03604_ _02671_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__mux2_1
X_05315_ net190 _01027_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__nor2_1
X_09083_ net208 _04329_ _04330_ net400 net919 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__a32o_1
X_06295_ net148 _01966_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10397__SET_B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ net451 net448 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__and3_1
X_05246_ _00957_ _00958_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05177_ _00888_ _00889_ _00873_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09985_ clknet_leaf_73_wb_clk_i _00090_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_122_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07066__B _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ net235 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
X_08867_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] _00941_ vssd1 vssd1
+ vccd1 vccd1 _04196_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07818_ _01058_ net172 vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ net314 _01450_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_8_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07749_ _01084_ net144 vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10760_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[7\]
+ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_09419_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] _04567_
+ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07810__A _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05463__A2_N _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10691_ clknet_leaf_34_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[23\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08117__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05984__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07212__A2 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10125_ clknet_leaf_43_wb_clk_i _00163_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10056_ clknet_leaf_61_wb_clk_i net756 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10368__RESET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05224__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10958_ net598 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_128_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06487__B1 _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10889_ net645 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_39_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08027__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06336__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06055__B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05100_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ _00817_ _00823_ net1022 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06080_ _00655_ _01766_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05031_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _00762_ vssd1
+ vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__nor2_1
Xhold128 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold139 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_78_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10874__549 vssd1 vssd1 vccd1 vccd1 _10874__549/HI net549 sky130_fd_sc_hd__conb_1
XFILLER_0_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] _04767_ _04790_
+ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__and3_1
X_06982_ _00714_ _02645_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__nor2_1
X_05933_ net271 _01625_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05118__C _00685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ _04071_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_1_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05864_ _01548_ _01550_ _01551_ _01555_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06714__A1 _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ _03063_ _03093_ _03072_ _02182_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08583_ _03621_ _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05795_ _01486_ _01487_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__nand2_4
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05134__B _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07534_ _02779_ _03092_ _01619_ _02119_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06478__B1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ net409 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net392 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout332_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__and2_1
X_06416_ _02087_ _02088_ _02089_ _01711_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07396_ _02990_ _02991_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06493__A3 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07690__A2 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09135_ _04321_ _04364_ _04365_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout120_X net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06347_ _02018_ _02020_ _02021_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09066_ _04307_ _04309_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06278_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] _01941_ _01948_ vssd1
+ vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05453__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ net1055 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_select
+ sky130_fd_sc_hd__and2b_1
X_05229_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] _00941_ vssd1 vssd1
+ vccd1 vccd1 _00942_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07077__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ clknet_leaf_83_wb_clk_i _00073_ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_51_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _04222_ _04223_ _04225_ _04227_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__or4b_2
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] _01777_
+ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07524__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06705__A1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10461__RESET_B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06181__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10812_ clknet_leaf_59_wb_clk_i _00633_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10743_ clknet_leaf_63_wb_clk_i _00573_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07130__A1 _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10674_ clknet_leaf_33_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[6\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07969__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05995__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__X _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07197__A1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07197__B2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05219__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ clknet_leaf_55_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\]
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10039_ _00059_ _00637_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06172__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05580_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01253_
+ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07250_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06201_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__inv_2
X_07181_ _02138_ net81 _02750_ _02831_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07449__X _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06132_ net125 _01699_ net156 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06063_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05014_ net263 net262 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07188__A1 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 net408 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_2
Xfanout416 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09822_ _04827_ _04834_ _04835_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__nor3_1
Xfanout427 net429 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_2
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout438 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\] vssd1 vssd1 vccd1
+ vccd1 net438 sky130_fd_sc_hd__clkbuf_2
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_1
X_09753_ _00652_ _04783_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__nor2_1
X_06965_ _02602_ _02634_ _02635_ _00746_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout282_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _01238_ _04062_ _01240_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__a21o_1
X_05916_ _01582_ _01597_ _01604_ net118 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__and4_2
XANTENNA__07344__B net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__inv_2
X_06896_ _02564_ _02565_ _02566_ _02486_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__or4b_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__B1 _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08635_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ _04062_ net455 vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__o21ai_1
X_05847_ _01508_ _01519_ _01539_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08566_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ _03614_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05778_ net410 _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__nor2_1
XANTENNA__05910__A2 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07517_ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07112__A1 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08497_ net53 net145 _03959_ net1073 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o31a_1
XANTENNA__08175__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07448_ team_07_WB.EN_VAL_REG net386 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__or2_1
XFILLER_0_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout89 _01606_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05674__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] _02979_
+ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ clknet_leaf_17_wb_clk_i net672 net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_09049_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ _04301_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__or2_1
XANTENNA__07966__A3 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06423__B _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold470 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold481 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net386 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
Xhold492 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ clknet_leaf_60_wb_clk_i _00556_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07654__A2 _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05996__Y _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10657_ clknet_leaf_19_wb_clk_i _00512_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload15 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_2
Xclkload26 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__bufinv_16
Xclkload37 clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_6
X_10588_ clknet_leaf_31_wb_clk_i _00452_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_sck
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload48 clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__clkinv_8
Xclkload59 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_114_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06668__A2_N _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07709__A3 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06750_ net173 _02418_ _02421_ _00971_ net137 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a221o_1
XANTENNA__08975__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05701_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] vssd1
+ vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__nor2_1
X_06681_ _02351_ _02353_ _02327_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08420_ net472 _03642_ _03665_ net465 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__o211ai_1
X_05632_ net440 _01327_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06696__A3 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05252__X _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08351_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] _03826_
+ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05563_ _01273_ _01275_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06508__B _02180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07302_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ _02925_ _02928_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[5\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08282_ _00717_ _03643_ net466 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05494_ _01204_ _01206_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10923__667 vssd1 vssd1 vccd1 vccd1 net667 _10923__667/LO sky130_fd_sc_hd__conb_1
XFILLER_0_116_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06227__C _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload9 clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_8
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07233_ net126 _02773_ _02883_ _02874_ _02767_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout128_A _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07164_ net107 _01710_ _02761_ _02781_ _02803_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_22_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06524__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06115_ net126 _01701_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08070__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07095_ _02109_ _02139_ _02735_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__o21a_1
XANTENNA__05959__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06243__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06046_ net124 _01700_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__nor2_2
Xfanout202 _04583_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
XFILLER_0_100_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout224 _04510_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
Xfanout246 _04729_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_2
XANTENNA_input2_A gpio_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _04823_ _04821_ net1026 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
Xfanout257 _01488_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_8
Xfanout268 _04591_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
X_07997_ _03548_ _03549_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__xnor2_1
Xfanout279 net281 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
XANTENNA__06384__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__and4_1
X_06948_ _02615_ _02616_ _02618_ _02614_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__or4b_1
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09667_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ _04721_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06879_ _02543_ _02529_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08618_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net455 vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09598_ _04666_ _04674_ _04676_ _04664_ net1043 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07090__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ net1145 _03610_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08914__A team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511_ clknet_leaf_12_wb_clk_i _00379_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ clknet_leaf_42_wb_clk_i _00326_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06434__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10373_ clknet_leaf_17_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[1\]
+ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05992__B net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06375__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06609__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__A2 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10709_ clknet_leaf_69_wb_clk_i _00540_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992__632 vssd1 vssd1 vccd1 vccd1 _10992__632/HI net632 sky130_fd_sc_hd__conb_1
XANTENNA__08052__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07920_ _03306_ _03445_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07851_ net161 _03366_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08760__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ net99 _02470_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__nand2_1
Xinput2 gpio_in[23] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_2
X_07782_ _01105_ _02212_ _02191_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__a21oi_1
X_04994_ net459 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
X_09521_ _00665_ _01419_ net289 _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__o211a_1
X_06733_ net420 net419 _02360_ _02361_ _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a311o_1
XFILLER_0_79_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10102__Q team_07_WB.instance_to_wrap.team_07.displayPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09452_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] net413
+ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o21ai_1
X_06664_ _01626_ _02258_ _01638_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _03858_ _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05615_ net442 net439 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__or2_1
X_09383_ net224 _04545_ _04546_ net395 net870 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06595_ net253 _02264_ _02265_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08334_ _03809_ _03810_ net488 vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05546_ net417 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01259_ sky130_fd_sc_hd__or3_2
XFILLER_0_129_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05710__X _01423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ net4 _00660_ _00663_ _03704_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a41o_1
X_05477_ _01153_ _01174_ _01189_ _01046_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__o22a_2
XFILLER_0_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08453__B _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07216_ _02065_ net82 _02736_ _02861_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ _00678_ net458 _01254_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07147_ net104 _02277_ _02761_ net164 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07078_ _02726_ _02729_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06029_ net134 net125 net144 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a21oi_4
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ _04754_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] vssd1 vssd1
+ vccd1 vccd1 _04760_ sky130_fd_sc_hd__a31o_1
X_10991_ net631 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06148__B _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06716__X _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05987__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10976__616 vssd1 vssd1 vccd1 vccd1 _10976__616/HI net616 sky130_fd_sc_hd__conb_1
XANTENNA__07490__B1 _03050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10425_ clknet_leaf_1_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[2\]
+ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10356_ clknet_leaf_56_wb_clk_i _00296_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10287_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[0\]
+ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08742__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06339__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05400_ _01056_ _01094_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06380_ _01662_ _01668_ _01663_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a21o_4
XFILLER_0_111_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05331_ _01035_ _01037_ _01043_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__or3b_1
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08050_ net1147 net295 _03578_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__a21o_1
X_05262_ _00673_ _00974_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07001_ _02664_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05193_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06802__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row net414 _04234_
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared vssd1 vssd1 vccd1
+ vccd1 _04243_ sky130_fd_sc_hd__a31o_1
XANTENNA__05726__C_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ net133 _03366_ _03365_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08328__A3 _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ _04206_ net436 _04205_ vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
XANTENNA__06240__C _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05137__B _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ net106 _03380_ _03388_ _01692_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07765_ _03319_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__inv_2
X_04977_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] vssd1
+ vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout362_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09504_ net934 net204 _04630_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06716_ net143 _01737_ _02260_ _02388_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07696_ _01619_ net249 _02249_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__or3b_1
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09435_ _01429_ _01430_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06647_ _02067_ _02281_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09366_ net224 _04532_ _04534_ net396 net1122 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a32o_1
X_06578_ net277 net98 net119 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08317_ _03742_ _03794_ _03793_ net484 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05529_ _01197_ _01240_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__nor2_1
X_09297_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _03725_ _03726_
+ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08179_ _03644_ _03656_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ clknet_leaf_72_wb_clk_i _00214_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06712__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect
+ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.flagPixel sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05786__B1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05328__A _01008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ clknet_leaf_62_wb_clk_i _00130_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07527__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05538__B1 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10974_ net614 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__06159__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05998__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08374__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06606__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05510__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07463__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10408_ clknet_leaf_18_wb_clk_i _00299_ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10339_ clknet_leaf_50_wb_clk_i _00279_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07230__A3 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07518__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05880_ _01569_ _01570_ _01572_ _01573_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__or4b_4
XFILLER_0_108_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08069__A_N net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07550_ net167 _02262_ _02219_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06501_ _02173_ _02174_ _02149_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07481_ _01658_ _01873_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09220_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06432_ net285 net282 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__or2_4
XFILLER_0_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06363_ net136 net125 net168 _01935_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06075__Y _01762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ _03603_ _03602_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05314_ _01010_ _01019_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__or2_1
X_09082_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a21o_1
X_06294_ net148 _01966_ _01969_ net160 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_114_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ _03568_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ net389 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__mux2_1
X_05245_ _00684_ _00946_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05176_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\]
+ _00883_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
X_09984_ clknet_leaf_72_wb_clk_i _00089_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ net235 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07066__C net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ _00685_ _04192_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07817_ _01058_ net172 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__nor2_1
X_08797_ net794 _04151_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07748_ _01068_ net157 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07679_ _03161_ _03234_ _03236_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__a21o_1
X_09418_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ _04572_ _04567_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
XANTENNA__07810__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10690_ clknet_leaf_34_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[22\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10667__RESET_B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09349_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06442__A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input40_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ clknet_leaf_44_wb_clk_i _00162_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10055_ clknet_leaf_62_wb_clk_i net764 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05999__Y _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ net597 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10888_ net644 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_26_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06336__B net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05571__C_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07987__B2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold107 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold118 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05030_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__or2_1
Xhold129 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[7\] vssd1 vssd1
+ vccd1 vccd1 net798 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08043__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06352__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06981_ _02645_ _02646_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__nor2_1
X_05932_ net271 _01625_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__and2_2
X_08720_ _04034_ _04082_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_47_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08651_ _04066_ _04071_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__and3_1
X_05863_ _01548_ _01550_ _01551_ _01555_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_1_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06714__A2 _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07602_ _03073_ _03160_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08582_ net1166 _03620_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nand2_1
X_05794_ _01486_ _01487_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07533_ _00759_ net99 _01607_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout158_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ net451 net409 vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__nor2_1
XANTENNA__07630__B _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06527__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09203_ net5 net1180 _04417_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
X_06415_ _01709_ _01720_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__nor2_1
X_07395_ net1110 _02988_ net477 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_33_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06246__B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06346_ net175 _02014_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__or2_4
XANTENNA__07427__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07978__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04313_ _04315_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__nor4_1
XFILLER_0_44_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06277_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] net256 _01951_ vssd1
+ vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout113_X net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08016_ net1013 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_right
+ sky130_fd_sc_hd__and2b_1
X_05228_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] net446 vssd1 vssd1
+ vccd1 vccd1 _00941_ sky130_fd_sc_hd__nand2_1
XANTENNA__06650__A1 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06650__B2 _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05159_ _00865_ _00866_ _00871_ _00858_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__a31o_1
XANTENNA__07077__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ clknet_leaf_80_wb_clk_i _00072_ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07805__B net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ _00724_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _00725_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_51_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ net842 net152 net150 _04886_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__a22o_1
XANTENNA__07093__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ net391 net389 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__o21a_1
XANTENNA__07524__C net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06705__A2 _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05700__A_N net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ clknet_leaf_59_wb_clk_i _00632_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06469__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10742_ clknet_leaf_62_wb_clk_i _00572_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06437__A _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07130__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10673_ clknet_leaf_33_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[5\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10430__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05995__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07197__A2 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06900__A _00746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ clknet_leaf_56_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10038_ _00058_ _00636_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841__516 vssd1 vssd1 vccd1 vccd1 _10841__516/HI net516 sky130_fd_sc_hd__conb_1
XFILLER_0_112_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06200_ _01863_ _01865_ _01864_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07409__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10100__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06131_ net130 net123 _01677_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__or3_4
XFILLER_0_83_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06062_ _00687_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01238_
+ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__or3b_1
XFILLER_0_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05013_ net262 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07188__A2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
X_09821_ _04825_ _04833_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a21oi_1
Xfanout417 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] vssd1
+ vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_2
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06810__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout439 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[2\] vssd1 vssd1 vccd1
+ vccd1 net439 sky130_fd_sc_hd__buf_2
XANTENNA__07184__Y _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\] _04777_ vssd1 vssd1
+ vccd1 vccd1 _04783_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06964_ _02487_ _02560_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__nand2_1
X_08703_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _04067_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__or2_1
X_05915_ _01582_ net118 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__and2_2
X_09683_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\] vssd1 vssd1 vccd1
+ vccd1 _04736_ sky130_fd_sc_hd__and3_1
X_06895_ net117 _02476_ _02528_ _02539_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout275_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05846_ _01519_ _01539_ _01508_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__o21ai_1
X_08634_ _01196_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__nand2_1
XANTENNA__07641__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08565_ _04012_ _04013_ _03996_ vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__o21a_1
X_05777_ _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07516_ _02108_ _02150_ _03071_ _03073_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08496_ net139 _03629_ _03960_ net811 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07112__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06856__D1 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ net899 _03021_ _03023_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[23\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07378_ _02979_ _02980_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09117_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06329_ net124 _01963_ _01965_ _01993_ _01641_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a41o_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09048_ _04301_ _04302_ net1169 net407 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__a2bb2o_1
Xhold460 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold471 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold482 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net387 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
Xhold493 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06387__B1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06926__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10725_ clknet_leaf_60_wb_clk_i _00555_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08382__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ clknet_leaf_19_wb_clk_i _00511_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_8
XANTENNA__08064__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ clknet_leaf_31_wb_clk_i _00451_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_sdi
+ sky130_fd_sc_hd__dfrtp_1
Xclkload27 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload38 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinv_8
Xclkload49 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_114_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07726__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05700_ net419 net420 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__nand2b_4
X_06680_ _00759_ _01627_ _02178_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05631_ _01319_ _01343_ _00680_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__and3b_1
X_08350_ _03637_ _03815_ _03766_ _03632_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05562_ _01266_ _01274_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ _02928_ _02929_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08281_ net465 _03756_ _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06302__B1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05493_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ _01205_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__xnor2_1
X_07232_ _01936_ _02873_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06853__B2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ _02059_ _02773_ _02775_ _02072_ _02815_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06524__B net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06114_ net171 net141 net184 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05408__A2 _01112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ _02737_ _02738_ _02740_ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06045_ net1141 _01633_ _01641_ _01730_ _01734_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ sky130_fd_sc_hd__a2111oi_2
Xclkbuf_leaf_62_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout203 _04583_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
XANTENNA__09555__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05708__X _01421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 _01503_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_4
Xfanout225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
XANTENNA_fanout392_A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
Xfanout247 _04270_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
X_09804_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] _04811_ _04818_
+ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__and3_1
Xfanout258 _00798_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_4
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_4
X_07996_ net450 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__xor2_1
XANTENNA__07581__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout180_X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06947_ net197 _02500_ _02509_ _02617_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] _04721_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a21oi_1
X_06878_ _02548_ _02546_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__nand2b_1
X_08617_ _04045_ net1150 _04044_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__mux2_1
X_05829_ _00712_ _01516_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09597_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06258__Y _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ net993 _03961_ _04002_ vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_46_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07097__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07097__B2 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08479_ _03926_ _03949_ _03950_ _03753_ _03751_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__o32a_1
XFILLER_0_108_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ clknet_leaf_12_wb_clk_i _00378_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ clknet_leaf_42_wb_clk_i _00325_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_135_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10372_ clknet_leaf_4_wb_clk_i net714 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05782__C_N _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout93_X net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07546__A _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[1\] vssd1 vssd1
+ vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06375__A3 _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06609__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07088__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07088__B2 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10708_ clknet_leaf_68_wb_clk_i _00539_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06625__A _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10639_ clknet_leaf_37_wb_clk_i _00503_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09936__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06360__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09001__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07850_ _01094_ net158 vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nor2_1
X_06801_ _01590_ _01598_ _02470_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__and3_1
X_07781_ _03281_ _03283_ _03299_ _03301_ _03276_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__o221a_1
X_04993_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1 vssd1
+ vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
Xinput3 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_2
X_09520_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _01420_
+ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand2_1
X_06732_ _02369_ _02378_ _02384_ _02404_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__or4b_1
XFILLER_0_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06663_ _02293_ _02294_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__or2_2
XANTENNA__05326__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ net961 net202 _04596_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10847__522 vssd1 vssd1 vccd1 vccd1 _10847__522/HI net522 sky130_fd_sc_hd__conb_1
XFILLER_0_8_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08402_ _00711_ _03876_ _03854_ _03718_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a211oi_1
X_05614_ net443 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1
+ vccd1 vccd1 _01327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09382_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04541_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__nand3_1
X_06594_ net255 _02265_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ team_07_WB.instance_to_wrap.team_07.circlePixel _03671_ net486 _00727_ vssd1
+ vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o211ai_2
X_05545_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout238_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08264_ _00663_ _03704_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05476_ net296 _01018_ _01182_ _01184_ _01188_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06535__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07215_ _01795_ _01901_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__and3_1
X_08195_ net486 _03673_ net488 vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06254__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07146_ _02793_ _02797_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07077_ net96 net89 net86 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__and3_2
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06028_ net169 _01715_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10934__583 vssd1 vssd1 vccd1 vccd1 _10934__583/HI net583 sky130_fd_sc_hd__conb_1
X_07979_ _03308_ _03441_ _03533_ _03496_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__o31a_1
X_09718_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] _04756_ _04757_
+ _04759_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__o22a_1
X_10990_ net630 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09649_ _00761_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05901__X _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06817__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05987__C _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06445__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10424_ clknet_leaf_1_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[1\]
+ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06045__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10355_ clknet_leaf_55_wb_clk_i _00295_ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09519__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ clknet_leaf_78_wb_clk_i _00278_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05067__Y _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__A1_N _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06339__B _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05330_ _01036_ _01041_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08046__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05261_ _00973_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07000_ _02662_ _02663_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05192_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00905_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07233__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07233__B2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07186__A _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ net491 _04242_ vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07902_ net257 _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__or2_1
X_08882_ _01966_ _04203_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07914__A _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _03381_ _03387_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _03311_ _03312_ _03318_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__nand3_2
X_10888__644 vssd1 vssd1 vccd1 vccd1 net644 _10888__644/LO sky130_fd_sc_hd__conb_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04976_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] vssd1
+ vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
X_09503_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ net268 _04627_ _04629_ net222 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__a221o_1
X_06715_ _01804_ _02044_ _02013_ net254 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__and4b_1
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ _02109_ net81 _02771_ _01637_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout355_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ _04556_ _03593_ _00813_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__mux2_2
XANTENNA__05153__B team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06646_ _02316_ _02317_ _02318_ _02313_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09365_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06577_ _02178_ _02249_ _02250_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] _03744_ _03780_
+ _03709_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a31o_1
X_05528_ _01238_ _01240_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__or2_1
X_09296_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04481_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08247_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\] _00730_ _03724_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] vssd1 vssd1 vccd1 vccd1
+ _03726_ sky130_fd_sc_hd__a31o_1
X_05459_ _01167_ _01168_ _01170_ _01171_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08178_ _00703_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nand2_2
XFILLER_0_127_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07224__A1 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07224__B2 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ _02277_ _02758_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06712__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect
+ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ clknet_leaf_46_wb_clk_i _00129_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07824__A _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__B1 _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10973_ net613 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05998__B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06175__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06606__C _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ clknet_leaf_18_wb_clk_i _00298_ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10338_ clknet_leaf_23_wb_clk_i net1161 net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10269_ clknet_leaf_8_wb_clk_i _00261_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07734__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08479__B1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06500_ _02139_ _02160_ _02166_ _02032_ _02159_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a221o_1
X_07480_ _01961_ _03038_ _03039_ _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_17_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06431_ _02062_ _02076_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a21o_1
XANTENNA__07900__C net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09150_ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__inv_2
X_06362_ net133 net128 _01935_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__and3_4
XFILLER_0_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08101_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__mux4_1
X_05313_ _01008_ _01025_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__nor2_1
X_09081_ _04328_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__inv_2
X_06293_ net437 _01968_ _01967_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08032_ net409 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net291 _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05244_ net456 _00956_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07909__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05175_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ _00883_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09983_ clknet_leaf_72_wb_clk_i _00088_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05148__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ net429 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XANTENNA__08299__X _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A2 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _04194_ _04193_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] vssd1
+ vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07816_ _03370_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__or3b_1
XFILLER_0_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08796_ _04151_ _04152_ net192 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_84_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07747_ _03299_ _03301_ _03286_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__nand3b_1
X_04959_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\] vssd1 vssd1
+ vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07678_ _03119_ _03153_ _03235_ _02697_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ _04570_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nor2_1
X_06629_ _02164_ _02301_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09348_ net223 _04519_ _04521_ net395 net864 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09279_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05456__B1 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__A _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06653__C1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06723__A _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ clknet_leaf_44_wb_clk_i _00161_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07554__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ clknet_leaf_62_wb_clk_i net767 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input33_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05345__Y _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08937__X _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10956_ net596 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__07133__B1 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06487__A2 _02042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10887_ net562 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XFILLER_0_39_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05080__Y _00807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold108 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold119 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06352__B _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09944__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06980_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _02643_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] vssd1 vssd1
+ vccd1 vccd1 _02646_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05931_ net283 _01623_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__nand2_4
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08650_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__xnor2_1
X_05862_ _01548_ _01555_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07601_ _03070_ _03093_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08581_ _04016_ _04024_ _03996_ vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__o21a_1
XANTENNA__10701__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05793_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] vssd1 vssd1
+ vccd1 vccd1 _01487_ sky130_fd_sc_hd__a41o_1
XFILLER_0_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07532_ _03084_ _03086_ _03090_ _03075_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06808__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05712__A _01424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ net391 net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ _03032_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[25\]
+ sky130_fd_sc_hd__a221o_1
XANTENNA__07675__A1 _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06527__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _04372_ _04413_ _04414_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__or4_1
X_06414_ _01675_ _01708_ net199 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__o21a_2
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07394_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\]
+ _02987_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__or4b_1
XFILLER_0_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06345_ _00710_ net131 _01698_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout318_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or4_1
X_06276_ net180 _01929_ _01948_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__o211a_1
XANTENNA__06543__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08015_ net1049 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_left
+ sky130_fd_sc_hd__and2b_1
X_05227_ _00883_ _00831_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_130_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06262__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout106_X net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05158_ _00867_ _00868_ _00869_ _00870_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__a22o_1
XANTENNA__07077__C net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05089_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__or2_1
X_09966_ clknet_leaf_82_wb_clk_i _00071_ net301 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_08917_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__xnor2_1
X_09897_ _01777_ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08848_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ net294 net291 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ _04184_ vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08779_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\] net399 net957
+ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10810_ clknet_leaf_67_wb_clk_i _00631_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06469__A2 _02101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07666__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ clknet_leaf_62_wb_clk_i _00571_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07130__A3 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ clknet_leaf_26_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[4\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05429__B1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07969__A2 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10470__RESET_B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05069__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07197__A3 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10106_ clknet_leaf_56_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\]
+ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10037_ _00057_ _00648_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08854__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sck vssd1 vssd1
+ vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09939__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10880__555 vssd1 vssd1 vccd1 vccd1 _10880__555/HI net555 sky130_fd_sc_hd__conb_1
XFILLER_0_26_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06130_ _01677_ _01692_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__nor2_2
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06363__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06061_ _00685_ _00828_ _00959_ _00961_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__or4_2
XFILLER_0_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10254__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05012_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] _00649_
+ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09820_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\] _04825_ _04833_
+ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__and3_1
Xfanout407 net408 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_2
Xfanout429 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] vssd1 vssd1 vccd1
+ vccd1 net429 sky130_fd_sc_hd__clkbuf_2
X_09751_ net244 _04780_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__nor2_1
X_06963_ _02479_ _02553_ _02633_ _02603_ _02557_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a311o_1
X_08702_ _01241_ _04112_ _04114_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__and3_1
X_05914_ _00716_ net128 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__xnor2_2
X_09682_ _04732_ _04733_ _04735_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__nor3_1
X_06894_ _02476_ _02528_ net117 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a21oi_1
X_08633_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__nand2_1
X_05845_ _01526_ _01529_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\]
+ _01523_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__o211a_1
XANTENNA__07896__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07641__B _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ net139 _03962_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__and2_1
XANTENNA__06538__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05776_ _01461_ _01467_ _01469_ _01474_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__nor4_4
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07515_ _02108_ _02150_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__o21a_1
XANTENNA__07648__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08495_ _03630_ _03961_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07446_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] _03021_
+ net230 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06320__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07377_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\] _02977_
+ _02974_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07369__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04347_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10228__RESET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06328_ _01985_ _01990_ _01999_ _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09047_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ _04299_ net248 vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06259_ net158 net146 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__nand2_8
XFILLER_0_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] vssd1 vssd1
+ vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\] vssd1 vssd1 vccd1
+ vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold472 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\] vssd1 vssd1
+ vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold483 team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06387__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09949_ net461 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05904__X _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10031__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10864__539 vssd1 vssd1 vccd1 vccd1 _10864__539/HI net539 sky130_fd_sc_hd__conb_1
XANTENNA__07639__A1 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06167__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724_ clknet_leaf_60_wb_clk_i _00554_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10655_ clknet_leaf_19_wb_clk_i _00510_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06454__Y _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload17 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__06183__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10586_ clknet_leaf_36_wb_clk_i _00450_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_ss
+ sky130_fd_sc_hd__dfstp_1
Xclkload28 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload39 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload39/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10206__Q team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05630_ _01331_ _01342_ _01337_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__or3b_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06358__A _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05561_ _01257_ _01264_ _01262_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07300_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08280_ _03637_ _03641_ _03657_ _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or4_1
X_05492_ net419 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07231_ _02033_ _02775_ _02872_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07162_ net104 _02277_ _02767_ net164 vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06113_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _00710_ _01436_
+ _01434_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] vssd1
+ vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a32o_1
X_07093_ _02152_ _02742_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06044_ net157 net124 _01732_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__o21ai_4
XANTENNA__06380__X _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout204 _04583_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_4
XANTENNA__06540__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 _04471_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
Xfanout237 net240 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09803_ _04821_ _04822_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__and2_1
Xfanout248 _04270_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_2
X_07995_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__xor2_1
Xfanout259 _00798_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
XANTENNA_fanout385_A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05156__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net1172 _04769_ _04770_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__a21bo_1
X_06946_ net211 _02510_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_31_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09665_ net1136 _04722_ _04723_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a21o_1
XANTENNA__07869__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06877_ net93 _02545_ _02547_ _02472_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout173_X net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _01929_ _01926_ _00964_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__mux2_1
X_05828_ _01509_ _01520_ _01507_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09596_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\]
+ _04672_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__and3_1
XANTENNA__06541__A1 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06268__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08547_ _03610_ _04001_ net140 vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a21o_1
X_05759_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08478_ net465 net470 _03664_ _03899_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o311a_1
XFILLER_0_64_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07429_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ _03008_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\] vssd1
+ vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_21_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10440_ clknet_leaf_42_wb_clk_i _00324_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10371_ clknet_leaf_3_wb_clk_i net688 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07827__A _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_07_WB.instance_to_wrap.ssdec_sdi vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06450__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout86_X net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08880__C_N net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__A _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06609__C _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ clknet_leaf_68_wb_clk_i _00538_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06625__B _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10638_ clknet_leaf_37_wb_clk_i _00502_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10569_ clknet_leaf_9_wb_clk_i _00437_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06599__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06360__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06800_ _02466_ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__nand2b_2
X_07780_ _03279_ _03334_ _03274_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06771__A1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04992_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel vssd1 vssd1
+ vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06771__B2 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06731_ _02386_ _02387_ _02392_ _02400_ _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06359__Y _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ net265 _04595_ net287 net217 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a221o_1
X_06662_ _01639_ _02259_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__nand2_1
X_10886__561 vssd1 vssd1 vccd1 vccd1 _10886__561/HI net561 sky130_fd_sc_hd__conb_1
XFILLER_0_59_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08401_ _03834_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__or2_1
X_05613_ net442 net441 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__and2_1
X_09381_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04538_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a31o_1
X_06593_ net253 _02021_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08332_ _03805_ _03808_ net485 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a21o_1
XANTENNA__08276__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05544_ net416 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01257_ sky130_fd_sc_hd__or3_2
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08263_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] _03741_
+ net487 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05475_ _01185_ _01186_ _01187_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout133_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06535__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07214_ _02134_ net82 _02741_ _02861_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08194_ net412 team_07_WB.instance_to_wrap.team_07.circlePixel _03672_ vssd1 vssd1
+ vccd1 vccd1 _03673_ sky130_fd_sc_hd__or3b_1
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07145_ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07076_ _02726_ _02729_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06027_ _01681_ _01716_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__or2_1
XANTENNA__07539__B1 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07978_ net132 _03304_ _03474_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ _00655_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] vssd1
+ vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06929_ _02588_ _02590_ _02598_ _02599_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_87_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09648_ _00655_ _04709_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_26_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _01793_ _03967_ _03976_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_65_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06285__X team_07_WB.instance_to_wrap.team_07.memGen.buttonHighlightDetect
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06445__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10423_ clknet_leaf_1_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[0\]
+ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ clknet_leaf_57_wb_clk_i _00294_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10285_ clknet_leaf_78_wb_clk_i _00277_ net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913__657 vssd1 vssd1 vccd1 vccd1 net657 _10913__657/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_109_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06505__A1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06636__A _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09947__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05260_ _00971_ _00972_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09758__A1 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05191_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ _00899_ _00900_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__mux4_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07233__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__S net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06371__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08950_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _00710_ _04234_
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared vssd1 vssd1 vccd1 vccd1
+ _04242_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07901_ _01058_ net214 _01723_ _03384_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__o22a_1
X_08881_ net437 _04205_ vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ _03382_ _03385_ _03386_ _03375_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__or4b_2
XFILLER_0_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07763_ _03317_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__inv_2
X_04975_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] vssd1
+ vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
X_09502_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\] vssd1
+ vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06714_ _02135_ _02259_ _02312_ _02140_ _02221_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__o221a_1
X_07694_ net112 _03249_ _01639_ _02760_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__or4b_1
X_09433_ _04557_ _03592_ _00813_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06645_ net282 _00757_ _02297_ _02308_ _02109_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout250_A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09364_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04530_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__and2_1
X_06576_ net93 net109 net96 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08315_ _03695_ _03792_ _03738_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05527_ _01239_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__nand2b_2
X_09295_ net225 _04483_ _04484_ net398 net1084 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08246_ _01284_ _01305_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05458_ _01002_ _01016_ _01035_ _01099_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ net469 _03655_ net465 vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__a21o_1
X_05389_ _00966_ _00967_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__or2_1
X_07128_ _02761_ _02764_ _02768_ _02781_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__a22o_1
XANTENNA__07224__A2 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06712__C _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07059_ _01630_ _02212_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10070_ clknet_leaf_48_wb_clk_i _00128_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07543__C net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06684__A_N _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972_ net612 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_104_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10982__622 vssd1 vssd1 vccd1 vccd1 _10982__622/HI net622 sky130_fd_sc_hd__conb_1
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07463__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ clknet_leaf_17_wb_clk_i net709 net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08412__A1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ clknet_leaf_25_wb_clk_i net679 net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_10268_ clknet_leaf_8_wb_clk_i _00260_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10199_ clknet_leaf_81_wb_clk_i _00203_ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__A1 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05934__C1 _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05822__X _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07151__B2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06430_ _02092_ _02103_ _02090_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08057__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06361_ net159 _01653_ _01685_ _01683_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__mux4_1
X_05312_ _00996_ _01010_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__or2_2
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09080_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06292_ net434 net436 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08031_ net452 net448 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05243_ _00953_ _00954_ _00955_ _00947_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__o31a_1
Xinput40 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05174_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00886_ vssd1 vssd1
+ vccd1 vccd1 _00887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06414__B1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08954__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ clknet_leaf_72_wb_clk_i _00087_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06965__B2 _00746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] net1160 net234 vssd1
+ vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06666__A2_N _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08864_ net446 net258 _04192_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__and3_1
X_07815_ _01057_ _01741_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__nor2_1
X_08795_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] _04147_ net948
+ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o21ai_1
X_10966__606 vssd1 vssd1 vccd1 vccd1 _10966__606/HI net606 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_84_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07746_ _03290_ _03300_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_84_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04958_ net1140 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ net199 _01723_ _01736_ _02829_ _03217_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _04568_ _04569_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06628_ _02296_ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09347_ _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06559_ _02228_ _02230_ _02232_ _02227_ _02226_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09278_ _04264_ net226 _04472_ net396 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06653__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08229_ net412 _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__nor2_1
XANTENNA__06282__Y _01959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07835__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ clknet_leaf_44_wb_clk_i _00160_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10034__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ clknet_leaf_61_wb_clk_i net839 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05355__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10955_ net595 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_86_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10886_ net561 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_38_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10209__Q team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold109 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10919__663 vssd1 vssd1 vccd1 vccd1 net663 _10919__663/LO sky130_fd_sc_hd__conb_1
XFILLER_0_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06947__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05930_ net284 net274 _01621_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07464__B net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05861_ _01538_ _01554_ _01542_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_1
X_07600_ _03069_ _03097_ _03125_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_1_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08580_ _03619_ _04023_ net140 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a21oi_1
X_05792_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__nand4_4
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07531_ _03081_ _03087_ _03089_ _02034_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__and4b_1
XFILLER_0_49_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07124__B2 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or4_1
X_06413_ net137 net105 net167 _02086_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a31o_2
XANTENNA__06527__C _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07393_ _02988_ _02989_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_33_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09132_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ _04327_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_33_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06344_ net414 net135 _02016_ _02018_ net127 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05438__A1 _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09063_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__or4b_1
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06275_ _01931_ _01949_ _01950_ _01951_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout213_A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ net1027 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_down
+ sky130_fd_sc_hd__and2b_1
X_05226_ _00685_ _00938_ _00828_ _00928_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__or4b_1
XFILLER_0_114_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08927__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05157_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00870_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05088_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__nor2_2
X_09965_ clknet_leaf_81_wb_clk_i _00070_ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_08916_ _00724_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _00725_ _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__a221o_1
X_09896_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] _01776_ vssd1
+ vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10016__RESET_B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ net392 net390 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08778_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ net399 vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__or3_2
XANTENNA__06558__X _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05462__X _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ _03277_ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07115__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10740_ clknet_leaf_62_wb_clk_i _00570_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07666__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10671_ clknet_leaf_33_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[3\]
+ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05069__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ clknet_leaf_48_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10036_ _00056_ _00647_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05904__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06909__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10938_ team_07_WB.instance_to_wrap.ssdec_sck vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10869_ net544 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_112_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06363__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06060_ _01457_ _01481_ _01483_ _00653_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05011_ _00635_ net285 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout408 _00807_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_4
Xfanout419 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[1\] vssd1
+ vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_4
X_09750_ _04767_ _04780_ _04781_ net244 net1164 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a32o_1
X_06962_ _02483_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__nand2_1
X_05913_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] net128
+ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__xnor2_2
X_08701_ _04120_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ _04115_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__mux2_1
X_09681_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ net246 vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__and3_1
X_06893_ net113 _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07345__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07345__B2 _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__nand2_1
XANTENNA__10699__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05844_ _01534_ _01537_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__nand2_1
XANTENNA__07922__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08563_ _03614_ _04011_ net139 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__a21oi_1
X_05775_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__or4b_1
XFILLER_0_77_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06538__B _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07514_ net100 _02191_ _03072_ _01612_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__o211ai_2
XANTENNA__07648__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ _03962_ net53 _03961_ vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ _03021_ _03022_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[22\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07376_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\] _02977_
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09115_ net209 _04352_ _04353_ net400 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06327_ _01987_ _01989_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06273__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ _00664_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_96_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06258_ net154 net144 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__nor2_2
XFILLER_0_60_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05209_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00922_ sky130_fd_sc_hd__nand2_1
Xhold440 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 net1109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06189_ net286 net134 _01848_ _01861_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold451 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] vssd1 vssd1 vccd1
+ vccd1 net1120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold473 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] vssd1 vssd1
+ vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _00201_ vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold495 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\] vssd1 vssd1 vccd1
+ vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06387__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07584__A1 _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09948_ net461 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ net833 net151 net149 _04874_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07324__S _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06448__B _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ clknet_leaf_57_wb_clk_i _00553_ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06847__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10654_ clknet_leaf_15_wb_clk_i _00509_ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06464__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08064__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ clknet_leaf_34_wb_clk_i _00449_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06183__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload18 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_4
Xclkload29 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_114_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10019_ clknet_leaf_33_wb_clk_i _00098_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05560_ _01270_ _01271_ _01269_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05491_ _01198_ _01200_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07230_ net126 net141 _02773_ _02877_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__a41o_1
XFILLER_0_129_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07161_ _02793_ _02798_ _02811_ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06112_ _00827_ _01789_ _01794_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a22o_1
XANTENNA__06524__D _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07092_ _01654_ net163 _01664_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a21o_1
XANTENNA__08460__C1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06043_ net155 net123 _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout205 _04583_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout216 _01502_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_8
Xfanout227 _04427_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
X_09802_ _04811_ _04818_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__a21o_1
Xfanout238 net240 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
Xfanout249 _02170_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
X_07994_ _03546_ _03547_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__xnor2_1
X_09733_ _00652_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] net244
+ _04768_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or4_1
X_06945_ net250 _02508_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout280_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] _04719_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 _04723_ sky130_fd_sc_hd__and4b_1
X_06876_ _01590_ _01598_ _02470_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a21oi_1
X_05827_ _01513_ _01516_ _00712_ _01507_ _01509_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a2111o_1
X_08615_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] _04044_ vssd1 vssd1
+ vccd1 vccd1 _00176_ sky130_fd_sc_hd__xnor2_1
X_09595_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] _04672_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_71_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08546_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ _03608_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__o21ai_1
X_05758_ _01454_ _01455_ _01456_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_46_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08477_ _03898_ _03948_ _03667_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05689_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\]
+ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\] team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\]
+ net438 net436 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07428_ net988 _03009_ _03011_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[16\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__06284__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06715__C _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] _02965_
+ _02967_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\] vssd1
+ vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_135_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10370_ clknet_leaf_3_wb_clk_i net699 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09029_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ _04286_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07827__B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold492_A team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _00099_ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
X_10831__506 vssd1 vssd1 vccd1 vccd1 _10831__506/HI net506 sky130_fd_sc_hd__conb_1
XANTENNA__05915__X _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06780__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950__590 vssd1 vssd1 vccd1 vccd1 _10950__590/HI net590 sky130_fd_sc_hd__conb_1
XANTENNA__07562__B _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06465__Y _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ clknet_leaf_68_wb_clk_i _00537_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10637_ clknet_leaf_37_wb_clk_i _00501_ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10568_ clknet_leaf_9_wb_clk_i _00436_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06599__A2 _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10499_ clknet_leaf_13_wb_clk_i _00367_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06641__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08745__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07548__B2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04991_ team_07_WB.instance_to_wrap.team_07.lcdOutput.stagePixel vssd1 vssd1 vccd1
+ vccd1 _00728_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput5 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06730_ _02402_ _02397_ _02394_ _02401_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06661_ _02108_ _02259_ _02333_ net89 net98 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__o221a_1
X_08400_ _03738_ _03871_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__o21a_1
X_05612_ net442 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__and2b_1
X_09380_ net224 _04543_ _04544_ net395 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__a32o_1
X_06592_ _02021_ _01654_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_47_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08331_ _00729_ _03736_ _03807_ _03738_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05543_ net416 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01256_ sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08262_ _00728_ _03740_ _03700_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__a21o_1
X_05474_ net426 net188 _01021_ _01062_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07213_ _02073_ _02862_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10542__RESET_B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08193_ team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel
+ team_07_WB.instance_to_wrap.team_07.flagPixel vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout126_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07144_ _02794_ _02796_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07075_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] net298 net297 team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\]
+ _02728_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06026_ net169 _01716_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07539__A1 _02080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07977_ net262 _03414_ _03416_ net263 vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _04757_ _04758_ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__and2_1
X_06928_ net131 _02497_ _02503_ _02596_ _02521_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_87_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _04703_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06859_ net117 _02471_ _02529_ net109 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__o22a_1
XANTENNA__06514__A2 _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07711__A1 _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09578_ _04637_ _04661_ net482 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_65_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ net1000 _03988_ vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_137_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06445__C net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10422_ clknet_leaf_18_wb_clk_i net235 net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_135_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07838__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10353_ clknet_leaf_57_wb_clk_i _00293_ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06461__B _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10284_ clknet_leaf_78_wb_clk_i _00276_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06202__A1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07950__A1 _03471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07702__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06636__B _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06269__B2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07748__A _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05190_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00901_ vssd1 vssd1
+ vccd1 vccd1 _00903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07610__A2_N _03144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08718__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07900_ _03384_ _03454_ net252 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__and3b_1
X_08880_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared _04204_ net487
+ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or3b_1
XFILLER_0_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07831_ _01094_ net183 vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__nor2_1
X_04974_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] vssd1
+ vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
X_07762_ _01076_ net187 _03316_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ net918 net204 _04628_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__o21a_1
X_06713_ _01732_ _02283_ _02385_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07693_ _00759_ net120 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__A1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ net1163 _04578_ _04579_ _04581_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__o22a_1
X_06644_ _02164_ _02295_ _02301_ _01921_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10723__RESET_B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04530_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__or2_1
X_06575_ _00754_ _02138_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08314_ _03791_ _01302_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__mux2_1
X_05526_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ _01196_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__and2_1
X_09294_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08245_ _01285_ _01306_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05457_ net432 _01072_ _01113_ _01036_ _01169_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout410_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08176_ net472 net470 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05388_ _01099_ _01100_ _01066_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07127_ _00755_ _01629_ _02780_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07058_ _01630_ _02209_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__nor2_1
XANTENNA__06712__D _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06009_ net134 net142 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09977__RESET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05906__A _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10971_ net611 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_134_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05912__Y _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07840__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07332__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05171__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07568__A _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10405_ clknet_leaf_17_wb_clk_i net672 net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10837__512 vssd1 vssd1 vccd1 vccd1 _10837__512/HI net512 sky130_fd_sc_hd__conb_1
XANTENNA__07620__B1 _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10336_ clknet_leaf_25_wb_clk_i net678 net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10267_ clknet_leaf_8_wb_clk_i _00259_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10198_ clknet_leaf_80_wb_clk_i _00202_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__A2 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05934__B1 _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07750__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06647__A _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07151__A2 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06366__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06360_ net130 net125 _01686_ _01936_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__or4_2
XANTENNA__05270__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05311_ net188 _01015_ _01023_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__o21ba_1
X_06291_ net434 _01397_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08030_ _03566_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net389 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05242_ net298 _00874_ _00900_ net297 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07478__A _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput41 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06382__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05173_ _00884_ _00885_ _00873_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_2
X_10894__650 vssd1 vssd1 vccd1 vccd1 net650 _10894__650/LO sky130_fd_sc_hd__conb_1
XANTENNA__06414__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07611__B1 _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ clknet_leaf_72_wb_clk_i _00086_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08932_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08863_ net446 _04192_ _04193_ vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__o21a_1
X_07814_ _01113_ net183 vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__nand2_1
X_08794_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\]
+ _04147_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__or3_1
XANTENNA__07941__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04957_ net7 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
X_07745_ _00753_ _03292_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout360_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07676_ _02040_ _02260_ _03198_ _01655_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09415_ net480 _02961_ _04556_ _00819_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o2bb2a_1
X_06627_ _02265_ _02294_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09346_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__and3_1
X_06558_ net122 net199 _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__o21a_2
XFILLER_0_48_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05509_ net420 net419 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__and2b_1
X_09277_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nand2_1
X_06489_ _02155_ _02162_ _02161_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08228_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03706_ vssd1
+ vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08159_ net472 _03640_ _03642_ _03638_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10121_ clknet_leaf_44_wb_clk_i _00159_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05907__Y _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07327__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ clknet_leaf_62_wb_clk_i _00110_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07851__A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input19_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ net594 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XANTENNA__07133__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10885_ net560 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_38_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06892__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10139__D team_07_WB.instance_to_wrap.team_07.recGen.circleDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06644__A1 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06644__B2 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ clknet_leaf_24_wb_clk_i net745 net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05546__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989__629 vssd1 vssd1 vccd1 vccd1 _10989__629/HI net629 sky130_fd_sc_hd__conb_1
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05860_ _01534_ _01536_ _01537_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05791_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] vssd1 vssd1
+ vccd1 vccd1 _01485_ sky130_fd_sc_hd__nand3_1
XANTENNA__06580__B1 _02230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07530_ net178 net169 _02082_ _02097_ _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__o311a_1
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07461_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net392 net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ _03031_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[24\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06332__B1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09200_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__or4b_1
X_06412_ net210 net138 _01706_ _02054_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_119_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07392_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] _02987_
+ net478 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ _04318_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_33_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06343_ _01724_ _02012_ _02017_ _02011_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__or4b_1
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06824__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06274_ _00684_ net456 net196 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05225_ _00935_ _00936_ _00937_ _00931_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__o31a_1
XFILLER_0_103_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08013_ net1042 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_up
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_25_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05156_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07936__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07060__A1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05087_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\]
+ _00812_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__or3_2
X_09964_ clknet_leaf_83_wb_clk_i _00069_ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08915_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__xor2_1
X_09895_ net841 net151 net149 _04884_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout196_X net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08846_ net741 _04183_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__and2_1
XANTENNA__06804__A1_N net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05374__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _04138_ net399 net1102 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
X_05989_ _01677_ _01679_ net169 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07390__B net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05903__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ _01065_ net118 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__nor2_1
XANTENNA__07115__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07659_ _01680_ net165 _02835_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__a21o_1
XANTENNA__08863__A2 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07666__A3 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ clknet_leaf_26_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[2\]
+ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09329_ _00662_ _04507_ _04508_ _04503_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08076__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06626__A1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07051__A1 _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ clknet_leaf_56_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\]
+ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_10035_ _00055_ _00646_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_19_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06909__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ team_07_WB.instance_to_wrap.ssdec_ss vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868_ net543 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__08616__S _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10770__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ clknet_leaf_70_wb_clk_i _00620_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06617__A1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05010_ team_07_WB.EN_VAL_REG net41 _00745_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06660__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout409 _00706_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06961_ _00695_ _02106_ _00749_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a21o_1
X_08700_ _04117_ _04118_ _04119_ net258 vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__o211a_1
X_05912_ _01596_ _01603_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__nor2_2
X_09680_ _00655_ _04703_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nand2_1
XANTENNA__06659__X _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06892_ net430 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _02466_ _02467_
+ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__o22a_1
X_08631_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__or3b_1
X_05843_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] _01520_
+ _01523_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__and3_1
X_08562_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ _03613_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06160__A1_N net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05774_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\] _01472_ vssd1
+ vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__or4b_1
XANTENNA__10233__SET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07513_ net94 net86 _02332_ net96 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ _03650_ _03652_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__nand2_1
XANTENNA__07648__A3 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout156_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07444_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\] _03019_
+ net481 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06835__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ _02977_ _02978_ _02974_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout323_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__nand2_1
X_06326_ net215 _01969_ _02000_ _02001_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09045_ net247 _04298_ _04300_ net407 net1052 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06257_ _01933_ _01925_ _01923_ _01932_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__nand4b_1
XTAP_TAPCELL_ROW_96_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05208_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00921_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold430 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\] vssd1
+ vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__dlygate4sd3_1
X_06188_ _01852_ _01868_ _01854_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a21oi_1
Xhold441 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\] vssd1 vssd1
+ vccd1 vccd1 net1110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07033__A1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05139_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00852_ sky130_fd_sc_hd__or2_1
Xhold474 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07385__B net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared vssd1 vssd1
+ vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06387__A3 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09947_ net461 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09878_ _01772_ _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__nand2_1
X_08829_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _04141_
+ net1056 vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10722_ clknet_leaf_67_wb_clk_i _00010_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05920__Y _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08049__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10018__SET_B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10653_ clknet_leaf_15_wb_clk_i _00508_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06464__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10584_ clknet_leaf_41_wb_clk_i _00448_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload19 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06480__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07024__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05824__A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ clknet_leaf_33_wb_clk_i _00097_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07348__A2_N team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05490_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01202_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07160_ _02058_ _02120_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06111_ _01789_ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ net250 _01657_ _01667_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__and3_1
X_06042_ net158 _01653_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__nand2_8
XFILLER_0_48_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout206 _04376_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
Xfanout217 net219 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
XFILLER_0_5_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09801_ _04811_ _04820_ _04808_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a21o_1
XANTENNA__05467__A_N _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 _04427_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_4
X_07993_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__xor2_1
X_09732_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] _04766_ _04769_
+ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__o21a_1
X_06944_ net182 _02612_ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__nor2_1
X_09663_ net1093 _04720_ _04722_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__o21a_1
XANTENNA__06526__B1 _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ net90 _02544_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__nand2_1
X_08614_ _04042_ _04043_ _00960_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a21o_1
X_05826_ _01513_ _01516_ _00712_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a21o_1
X_09594_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] _04664_ _04666_
+ _04673_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ _03609_ _04000_ _03999_ vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a21oi_1
X_05757_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _01453_ vssd1 vssd1
+ vccd1 vccd1 _01456_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _03755_ _03819_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05688_ _00681_ net436 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_98_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07427_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] _03009_
+ net230 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_40_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_21_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07358_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\]
+ _02966_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__or4b_1
XFILLER_0_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06057__A2 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06309_ net171 _01973_ _01984_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07289_ net440 _01326_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__nor2_1
X_09028_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ _04286_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold260 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\] vssd1 vssd1
+ vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05347__C _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870__545 vssd1 vssd1 vccd1 vccd1 _10870__545/HI net545 sky130_fd_sc_hd__conb_1
XANTENNA__07335__S _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06475__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10705_ clknet_leaf_68_wb_clk_i _00536_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07493__A1 _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10636_ clknet_leaf_37_wb_clk_i net896 net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10567_ clknet_leaf_10_wb_clk_i _00435_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10498_ clknet_leaf_14_wb_clk_i _00366_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06360__D _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07753__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04990_ net412 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
Xinput6 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_X clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06660_ net278 _01609_ _02031_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__and3_1
XANTENNA__07181__B1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05611_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] net440
+ team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] _01323_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__o32a_1
XFILLER_0_8_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06591_ net123 _01654_ _02261_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__or3_2
XANTENNA__05731__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08330_ net457 _03734_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05542_ net415 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] vssd1 vssd1 vccd1
+ vccd1 _01255_ sky130_fd_sc_hd__or3_2
XANTENNA__06385__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07484__A1 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ team_07_WB.instance_to_wrap.team_07.buttonPixel team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05473_ _01036_ _01037_ _01106_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07212_ _01653_ _01665_ net184 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_41_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08192_ team_07_WB.instance_to_wrap.team_07.flagPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel
+ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_41_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07143_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] net299 net394 _02795_
+ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06391__Y _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\] net299 net394 _02727_
+ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XANTENNA__05729__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06025_ net215 net195 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__nand2_1
X_10854__529 vssd1 vssd1 vccd1 vccd1 _10854__529/HI net529 sky130_fd_sc_hd__conb_1
XANTENNA__07539__A2 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07976_ _03280_ _03522_ _03530_ _03515_ _03518_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__o2111a_1
X_09715_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] net246 _04752_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\] vssd1 vssd1 vccd1
+ vccd1 _04758_ sky130_fd_sc_hd__a31o_1
X_06927_ _02593_ _02594_ _02596_ _02597_ _02589_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09646_ _01767_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06858_ net430 _02528_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__nand2_1
X_05809_ _01494_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__or3_1
X_09577_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] _04661_
+ _04663_ _04640_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _02410_ _02415_ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_26_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08528_ net1118 _03987_ vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_137_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06295__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08459_ _03714_ _03749_ _03751_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08941__C _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__A1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ clknet_leaf_56_wb_clk_i _00312_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07227__B2 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ clknet_leaf_57_wb_clk_i _00292_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05789__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10283_ clknet_leaf_79_wb_clk_i _00275_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05926__X _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07163__B1 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06476__Y _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06269__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07218__A1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ clknet_leaf_37_wb_clk_i _00483_ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07748__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10957__597 vssd1 vssd1 vccd1 vccd1 _10957__597/HI net597 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06729__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ _03383_ _03384_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__or2_1
XANTENNA__05284__A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ _03314_ _03315_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__nand2b_1
X_04973_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] vssd1
+ vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
X_09500_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ net268 _04625_ _04627_ net222 vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a221o_1
X_06712_ net250 _01734_ _02021_ _02154_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__or4_1
X_07692_ _03041_ _03247_ _03248_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recMOD.modSquaresDetect
+ sky130_fd_sc_hd__o21ba_1
X_09431_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ _04569_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06643_ _02031_ _02281_ _02314_ _02315_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_91_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06827__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ net223 _04529_ _04531_ net398 net1060 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__a32o_1
X_06574_ _02075_ _02098_ _02247_ net249 net87 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__o311a_1
XFILLER_0_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08313_ _01381_ _03733_ _03789_ _03790_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_129_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05525_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01237_ _01236_ _01234_ _01194_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a2111oi_4
X_09293_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout236_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08244_ net484 net412 _03721_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05456_ _01006_ _01056_ _01063_ _01058_ _01052_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06843__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08175_ _00733_ net129 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout403_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05387_ net188 _01014_ _01021_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__nor3_1
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06562__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07126_ net281 _00749_ _01607_ _01634_ _02779_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a311o_1
XFILLER_0_42_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07057_ _01811_ _02036_ _02709_ _02711_ _01903_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_58_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06008_ net130 _01698_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05906__B _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07959_ _00970_ _01058_ net115 _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a31o_1
XANTENNA__05943__A1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ net610 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
X_09629_ net984 _04696_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__xor2_1
XANTENNA__06499__A2 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06737__B net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05360__C _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08951__A_N net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07568__B _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08948__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ clknet_leaf_16_wb_clk_i net707 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10876__551 vssd1 vssd1 vccd1 vccd1 _10876__551/HI net551 sky130_fd_sc_hd__conb_1
XANTENNA__07620__A1 _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10335_ clknet_leaf_25_wb_clk_i net674 net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10266_ clknet_leaf_7_wb_clk_i _00258_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10197_ clknet_leaf_82_wb_clk_i net1153 net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__A3 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05934__A1 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07590__Y _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07151__A3 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05310_ net189 _01010_ _01021_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__nor3_2
X_06290_ _01397_ _01399_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05241_ net447 _00843_ net394 _00832_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__a31o_1
Xinput20 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10174__RESET_B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput31 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_1
XFILLER_0_71_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10257__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05172_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\]
+ _00883_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07611__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06414__A2 _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ clknet_leaf_81_wb_clk_i _00085_ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ net430 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XANTENNA__04911__A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ net446 net232 _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06178__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _01112_ net187 _01658_ _01057_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__a22o_1
X_08793_ _04149_ _04150_ net192 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07744_ _01064_ net108 _03280_ _03284_ _01609_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_84_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04956_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1 vccd1
+ vccd1 _00696_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06838__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _03162_ _03226_ _03232_ _03076_ _03225_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__a221o_1
XANTENNA__07678__B2 _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout353_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09414_ net480 _02961_ _04557_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06626_ _02109_ _02295_ _02297_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_47_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09345_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04514_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06557_ _01654_ _01829_ _01661_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07669__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05508_ _00691_ _01198_ _01203_ _00692_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a22o_1
X_09276_ net226 net396 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__mux2_1
X_06488_ _01655_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08227_ net2 _03704_ _03705_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__a31o_1
X_05439_ _01151_ _01126_ _00965_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _03640_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07109_ _01694_ net162 _02758_ _02761_ _02762_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ _03597_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ net229 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05917__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_A _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ clknet_leaf_44_wb_clk_i _00158_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10051_ clknet_leaf_62_wb_clk_i _00109_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06748__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10953_ net593 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10884_ net559 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_14_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07624__A2_N _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08397__A2 _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07585__Y _03144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10318_ clknet_leaf_24_wb_clk_i net802 net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ clknet_leaf_74_wb_clk_i _00241_ net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07109__B1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05790_ net1086 _00797_ _00827_ net483 vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a22o_1
XANTENNA__06580__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07460_ net453 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__and2b_1
XANTENNA__06332__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06411_ net137 net105 net167 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__and3_1
XANTENNA__10355__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07391_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] _02987_
+ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09130_ net400 _04324_ _04363_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06342_ _00710_ net216 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09061_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04309_ _04311_ _04307_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06273_ net456 net212 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ _03558_ _03559_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__xnor2_1
X_05224_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00937_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07495__Y _03055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05155_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00868_ sky130_fd_sc_hd__nand2_1
X_10972__612 vssd1 vssd1 vccd1 vccd1 _10972__612/HI net612 sky130_fd_sc_hd__conb_1
XANTENNA_fanout101_A _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05086_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ clknet_leaf_81_wb_clk_i _00068_ net301 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_65_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__xor2_1
XANTENNA__04998__D net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ _01776_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07952__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _04182_ _04183_ _04144_ vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06020__B1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_X net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ net399 _01457_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__nor2_1
XANTENNA__06571__A1 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05988_ net185 net177 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__or2_2
X_07727_ _01064_ net115 _03281_ _03276_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__o31a_1
XANTENNA__08848__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04939_ net440 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XANTENNA__06287__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ _01902_ _02087_ _03213_ _03215_ _03119_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06609_ net160 net125 _01652_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__and3_2
XFILLER_0_137_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07589_ net251 _03146_ _03147_ _03145_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a31o_1
X_09328_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ net397 _04259_ net225 vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__a22o_1
XANTENNA__09273__A0 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06087__B1 _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ _04458_ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07338__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07051__A2 _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ clknet_leaf_61_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\]
+ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_8_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input31_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _00054_ _00645_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_19_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10936_ team_07_WB.instance_to_wrap.ssdec_sdi vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07511__B1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10867_ net542 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05716__A_N net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ clknet_leaf_70_wb_clk_i _00619_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07102__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06363__D _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06660__B _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06005__X _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06960_ _02602_ _02604_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a21oi_1
X_05911_ _01597_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__nand2_1
XANTENNA__08220__X _03699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06891_ _02556_ _02561_ _02543_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a21o_1
X_08630_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04046_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__a31o_1
X_05842_ _01527_ _01535_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06388__A _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05292__A _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ net139 _04010_ _03963_ vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05773_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__and4b_1
X_07512_ _01628_ _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06675__X _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ net993 _03961_ vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07443_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ _03018_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07374_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a31o_1
XANTENNA__09211__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09113_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06325_ net256 _01397_ net434 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__or3b_1
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09044_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__inv_2
X_06256_ _00684_ net176 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_96_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10822__497 vssd1 vssd1 vccd1 vccd1 _10822__497/HI net497 sky130_fd_sc_hd__conb_1
X_05207_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00920_ sky130_fd_sc_hd__or2_1
Xhold420 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\] vssd1 vssd1
+ vccd1 vccd1 net1089 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout104_X net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06187_ _01855_ _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__nor2_1
Xhold431 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold442 team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] vssd1 vssd1 vccd1
+ vccd1 net1111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
X_05138_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00851_ sky130_fd_sc_hd__or2_1
Xhold464 team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\] vssd1 vssd1 vccd1
+ vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold486 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09946_ net463 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
X_05069_ net491 _00796_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06792__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\] vssd1 vssd1 vccd1
+ vccd1 _04873_ sky130_fd_sc_hd__o21ai_1
XANTENNA__05914__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\]
+ _04141_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__or3_1
XANTENNA__06544__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06298__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08759_ net953 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05930__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ clknet_leaf_56_wb_clk_i _00552_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08049__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10652_ clknet_leaf_15_wb_clk_i _00507_ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10583_ clknet_leaf_41_wb_clk_i _00447_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06480__B net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05377__A _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ clknet_leaf_31_wb_clk_i _00096_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05824__B _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06001__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10919_ net663 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06110_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\] _01792_ vssd1 vssd1
+ vccd1 vccd1 _01793_ sky130_fd_sc_hd__and4b_2
XFILLER_0_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07090_ net251 _01657_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__nand2_2
XANTENNA__08460__A1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06671__A _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06041_ net156 _01652_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07486__B _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05287__A _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout207 _04376_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
X_09800_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] _04818_ vssd1
+ vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nand2_1
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_2
Xfanout229 _03594_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07992_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ net1134 vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__xor2_1
X_09731_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _04768_ net244
+ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a21o_1
X_06943_ net182 _02612_ _02613_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a21oi_1
X_09662_ _04716_ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor2_1
X_06874_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__inv_2
XANTENNA__06526__A1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__B1 _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _00964_ _01927_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nand2_1
X_05825_ _00712_ net196 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09593_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] _04672_ vssd1
+ vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08544_ net849 _03608_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__nand2_1
X_05756_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] vssd1 vssd1 vccd1
+ vccd1 _01455_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_46_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08475_ _03908_ _03946_ net489 _03753_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_46_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05687_ _00681_ net436 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07426_ _03009_ _03010_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[15\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07357_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06308_ _00681_ net180 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__nand2_1
XANTENNA__06057__A3 _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07288_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09027_ net247 _04285_ _04287_ net404 net859 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06239_ net101 _01825_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold250 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold272 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] vssd1 vssd1
+ vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout81_A _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05925__A _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10458__RESET_B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _00701_ _01786_ net152 _04904_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__o31a_1
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05931__Y _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06756__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10704_ clknet_leaf_68_wb_clk_i _00535_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07493__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10635_ clknet_leaf_38_wb_clk_i _00499_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10566_ clknet_leaf_6_wb_clk_i _00434_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06491__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10497_ clknet_leaf_13_wb_clk_i _00365_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07462__A_N net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06205__B1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__Y _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput7 wb_rst_i vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07181__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05610_ net442 net441 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__or2_1
X_06590_ net123 _01654_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__or2_1
XANTENNA__05731__A2 _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05541_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] vssd1 vssd1 vccd1
+ vccd1 _01254_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06385__B _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _03737_ _03738_ net485 vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05472_ _01059_ _01088_ _01068_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07211_ _02138_ net82 _02750_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08191_ _03658_ _03666_ _03669_ _03630_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07142_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\]
+ net446 vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06444__B1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07073_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\]
+ net446 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05729__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06024_ net195 net201 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__nand2_2
XFILLER_0_112_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07975_ _03346_ _03432_ _03528_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09714_ _04733_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__nor2_1
X_06926_ net428 net148 _02581_ _02501_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _04705_ _04706_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__or4_2
X_06857_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout171_X net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05808_ _01494_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__nor3_1
X_09576_ _04637_ _04661_ net482 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__o21ai_1
X_06788_ _01626_ _02412_ _02459_ _01636_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05480__A _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] _03980_ _03985_
+ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05739_ net1128 _00791_ _01441_ _00766_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _03877_ _03930_ net490 net462 _03858_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_19_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07409_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] _02998_
+ net230 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] vssd1 vssd1 vccd1
+ vccd1 _03864_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ clknet_leaf_56_wb_clk_i _00311_ net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05479__X _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10351_ clknet_leaf_33_wb_clk_i _00291_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10282_ clknet_leaf_73_wb_clk_i _00274_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout84_X net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09561__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05390__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06674__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10618_ clknet_leaf_38_wb_clk_i _00482_ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07218__A2 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07110__A _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06426__B1 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10549_ clknet_leaf_11_wb_clk_i _00417_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10244__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06729__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__B2 _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__B1 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06013__X team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07760_ _01067_ net216 net198 _01078_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__o22a_1
XANTENNA__05284__B net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04972_ net488 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
X_06711_ _02260_ _02262_ _02379_ _02383_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07691_ _01726_ _02365_ _03150_ _01712_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o22a_1
X_09430_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ _04577_ _04580_ _04568_ _04579_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__o221a_1
X_06642_ _02108_ _02209_ _02289_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06396__A _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04909__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__inv_2
X_06573_ _01687_ _01690_ _02049_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08312_ _00731_ _01303_ _03677_ _00732_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_19_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_05524_ _01220_ _01232_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__nand2_1
X_09292_ net226 _04480_ _04482_ net396 net889 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07457__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08243_ net484 net412 _03721_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05455_ _01156_ _01157_ _01158_ _01159_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout131_A _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ _03628_ _03648_ _03634_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05386_ net191 _01000_ _01021_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__nor3_2
XFILLER_0_70_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06417__B1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ net99 _01616_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07056_ _02688_ _02710_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__nor2_1
X_06007_ net144 net133 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_58_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07958_ _03509_ _03511_ _03512_ _03461_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a211o_1
XANTENNA__05943__A2 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] net160 vssd1 vssd1
+ vccd1 vccd1 _02580_ sky130_fd_sc_hd__nand2_1
X_07889_ _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09628_ _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_104_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06353__C1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ net828 net241 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07689__X team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06120__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06753__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10403_ clknet_leaf_17_wb_clk_i net680 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08948__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09556__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ clknet_leaf_26_wb_clk_i net700 net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07620__A2 _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10265_ clknet_leaf_7_wb_clk_i _00257_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10196_ clknet_leaf_80_wb_clk_i _00200_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05934__A2 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout390 _03562_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06344__C1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07105__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06944__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07111__Y _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05240_ net299 _00951_ _00952_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput43 wbs_we_i vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
X_05171_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\]
+ _00883_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07611__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ net432 net818 net236 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08861_ net240 _04191_ _01748_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__o21a_2
XANTENNA__06178__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ _03365_ _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__or2_1
X_08792_ net1015 _04147_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__nand2_1
X_07743_ _03282_ _03287_ _03295_ _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__a22o_1
X_04955_ net430 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XANTENNA__07127__A1 _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout179_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07674_ _02055_ _02282_ _03227_ _03231_ _01690_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a2111o_1
X_09413_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _02965_ _04557_ _02964_
+ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a2bb2o_1
X_06625_ _02031_ _02119_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09344_ net223 _04517_ _04518_ net399 net1057 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__a32o_1
X_06556_ _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05507_ _01219_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
X_09275_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ net1 net322 _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o211a_1
XANTENNA__07669__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06487_ _02039_ _02042_ _02152_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08226_ net4 net3 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nor2_1
X_05438_ _00966_ _00969_ _01136_ _01150_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08157_ net468 net470 vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05369_ _01079_ _01081_ _01078_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ net155 _01688_ net162 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08088_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ _00814_ net476 vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07039_ _02164_ _02362_ _02184_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05917__B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10050_ clknet_leaf_62_wb_clk_i _00108_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06574__C1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05933__A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10952_ net592 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_74_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10883_ net558 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06764__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10317_ clknet_leaf_24_wb_clk_i net834 net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_10248_ clknet_leaf_74_wb_clk_i _00240_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06004__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05546__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10179_ clknet_leaf_20_wb_clk_i _00189_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07109__A1 _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06332__A2 _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06410_ _02052_ _02083_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__nand2_1
X_07390_ _02987_ net478 _02986_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06341_ _01649_ _02011_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_33_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06393__B _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04310_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o21a_1
X_06272_ _00684_ net456 net196 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08011_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05223_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00936_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10324__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07045__B1 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05154_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00867_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07596__A1 _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05085_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00810_ vssd1 vssd1 vccd1
+ vccd1 _00811_ sky130_fd_sc_hd__nand2_1
X_09962_ clknet_leaf_79_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[39\]
+ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08913_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__xor2_1
X_09893_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] _01775_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ _04143_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_51_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06849__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06020__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05987_ net132 net128 _01676_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__and3_2
X_08775_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] net695 net238 vssd1
+ vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout463_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ net108 _03280_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04938_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] vssd1
+ vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout251_X net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ _03204_ _03214_ _03205_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a21oi_1
X_10827__502 vssd1 vssd1 vccd1 vccd1 _10827__502/HI net502 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06608_ _02268_ _02272_ _02273_ _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o22a_1
X_07588_ _01739_ _03078_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ net225 _04506_ _04507_ net396 net905 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a32o_1
X_06539_ net120 _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__or2_1
XANTENNA__08076__A2 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09258_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ _04454_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08209_ net417 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1 vssd1 vccd1 vccd1
+ _03688_ sky130_fd_sc_hd__and3b_1
X_09189_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10102_ clknet_3_0_0_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.displayDetect
+ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.displayPixel
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ _00053_ _00644_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06759__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06011__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__D1 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10935_ net584 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_105_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07511__A1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866_ net541 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ clknet_leaf_70_wb_clk_i _00618_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10995__635 vssd1 vssd1 vccd1 vccd1 _10995__635/HI net635 sky130_fd_sc_hd__conb_1
XFILLER_0_34_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07578__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06660__C _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05910_ _01583_ net121 _01602_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a21o_1
X_06890_ _02482_ _02560_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__nand2_1
X_05841_ _01524_ _01525_ _01529_ _01522_ _01521_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a32o_1
X_08560_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ _03613_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__xor2_1
X_05772_ _01463_ _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07511_ net89 net88 _01626_ net98 vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08491_ net139 _03960_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07442_ _03019_ _03020_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[21\]
+ sky130_fd_sc_hd__nor2_1
X_07373_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ _02969_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09112_ net209 _04349_ _04351_ net400 net1080 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06324_ net434 _01396_ _01489_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06255_ net212 _01926_ _01929_ net194 _01930_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout211_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05206_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold410 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] vssd1 vssd1
+ vccd1 vccd1 net1079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06186_ _01856_ _01857_ _01863_ _01866_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o22a_1
Xhold421 _04697_ vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] vssd1 vssd1
+ vccd1 vccd1 net1112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05137_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00850_ sky130_fd_sc_hd__nand2_1
Xhold454 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\] vssd1 vssd1
+ vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold476 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold498 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] vssd1 vssd1 vccd1
+ vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ net461 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
X_05068_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back _00795_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select vssd1
+ vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_5_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ net913 _04871_ _04872_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__o21a_1
X_08827_ _04171_ _04172_ net193 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07741__A1 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08758_ net997 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07709_ net155 net200 net170 _01744_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08689_ _00707_ _04105_ _04108_ _04110_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__o31a_1
XFILLER_0_135_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05930__B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ clknet_leaf_57_wb_clk_i _00551_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_fl_enable
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.sck_fl_enable
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10246__RESET_B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10979__619 vssd1 vssd1 vccd1 vccd1 _10979__619/HI net619 sky130_fd_sc_hd__conb_1
XFILLER_0_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ clknet_leaf_41_wb_clk_i _00446_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08733__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07980__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ clknet_leaf_31_wb_clk_i net898 net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06639__D net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06001__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10918_ net662 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10849_ net524 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XFILLER_0_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08445__C1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06952__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07767__B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06671__B _02027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06040_ net170 _01715_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06016__X _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout208 _04325_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
Xfanout219 _04582_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_1
XFILLER_0_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07991_ net257 _03437_ _03450_ _03505_ _03545_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recGen.circleDetect
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09730_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__nand2_1
X_06942_ _02500_ _02509_ net197 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06399__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05982__B1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] _04720_ vssd1
+ vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__and2_1
X_06873_ _02466_ _02474_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__or2_1
XANTENNA__06526__A2 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ _01109_ _01926_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand2_1
X_05824_ _01513_ _01516_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__nand2_1
X_09592_ _04665_ _04672_ _04669_ net1076 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_55_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10757__RESET_B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08543_ _03608_ _03995_ _03999_ vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__a21oi_1
X_05755_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\] vssd1 vssd1 vccd1
+ vccd1 _01454_ sky130_fd_sc_hd__or3_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05686_ net437 net436 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__or2_1
X_08474_ _03911_ _03930_ _03945_ net411 vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07425_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] _03008_
+ net478 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07356_ net482 _02963_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_21_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06307_ net184 _01975_ _01982_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_135_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07287_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09026_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06462__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06238_ _01888_ _01910_ _01916_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06169_ _01849_ _01809_ _01817_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__and3b_1
Xhold240 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] vssd1 vssd1
+ vccd1 vccd1 net909 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\] vssd1 vssd1
+ vccd1 vccd1 net942 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07693__A _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\] vssd1 vssd1 vccd1
+ vccd1 net953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] vssd1 vssd1
+ vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09928_ net341 _01785_ _01790_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a31o_1
X_09859_ _04666_ _04731_ _04767_ net264 team_07_WB.instance_to_wrap.audio vssd1 vssd1
+ vccd1 vccd1 _04861_ sky130_fd_sc_hd__o41a_1
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05941__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10703_ clknet_leaf_67_wb_clk_i _00534_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05899__B1_N _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09559__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ clknet_leaf_38_wb_clk_i net854 net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10565_ clknet_leaf_6_wb_clk_i _00433_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06491__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10496_ clknet_leaf_14_wb_clk_i _00364_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07108__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08902__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05540_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07469__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06385__C net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05471_ _01034_ _01080_ _01183_ _01145_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__o31a_1
XFILLER_0_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07210_ _02856_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__or2_1
X_08190_ _03631_ _03668_ _00717_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__mux2_1
XANTENNA__06682__A _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07141_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] net298 net297 team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05298__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07072_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] net298 _00942_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\]
+ _02725_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06023_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\] _01633_ _01641_
+ _01713_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_113_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07974_ _03340_ _03425_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07018__A team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\] net246 _04754_
+ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__and3_1
X_06925_ _02593_ _02595_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__nor2_1
X_09644_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__or4b_1
X_06856_ _02475_ _02492_ _02493_ _02526_ _01689_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05807_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nor2_2
X_09575_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] _04661_
+ _04662_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout164_X net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06787_ _00674_ _02332_ _02170_ net426 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a211oi_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _03980_ _03985_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__nand2_1
XANTENNA__05480__B _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05738_ _00652_ _00773_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08457_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03744_ _03804_
+ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__or4_2
XANTENNA__06132__B1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05669_ _01381_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07408_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] _02998_
+ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__and2_1
XANTENNA__07880__B1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08388_ net780 _03653_ _03832_ _03863_ vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07339_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _02411_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__A3 _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10350_ clknet_leaf_33_wb_clk_i _00290_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_115_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__and4_1
XFILLER_0_130_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10281_ clknet_leaf_82_wb_clk_i _00273_ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05936__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08031__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05942__Y _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07163__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06123__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06674__A1 _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10617_ clknet_leaf_40_wb_clk_i _00481_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07110__B _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07623__B1 _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ clknet_leaf_11_wb_clk_i _00416_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06007__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10479_ clknet_leaf_28_wb_clk_i _00347_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06729__A2 _02149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04971_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col vssd1 vssd1 vccd1
+ vccd1 _00710_ sky130_fd_sc_hd__inv_2
XANTENNA__08876__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06710_ _02154_ _02260_ _02382_ _02381_ _02380_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a32o_1
X_07690_ _01631_ _02009_ _02348_ net94 net100 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06641_ _00635_ _02212_ _02305_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_86_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06396__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09360_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__and3_1
X_06572_ net199 _02066_ _02171_ _02164_ _02158_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ net460 _01308_ _01384_ _03788_ net459 vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a311o_1
X_05523_ _01220_ _01232_ _01235_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__o22a_1
X_09291_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__inv_2
XANTENNA__06114__B1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08242_ _03672_ _03720_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__nor2_1
X_05454_ net296 _01029_ _01092_ _01154_ _01155_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__a221o_1
X_10860__535 vssd1 vssd1 vccd1 vccd1 _10860__535/HI net535 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_60_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06665__B2 _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_59_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_132_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08173_ _03628_ _03648_ _03634_ vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__a21o_1
X_05385_ _01096_ _01097_ _01094_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_132_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout124_A _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06417__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ _02729_ _02763_ _02777_ _01646_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07055_ _02681_ _02677_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06006_ net148 net131 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nor2_4
XFILLER_0_88_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07917__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__B2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _03288_ _03391_ _03351_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] net160 vssd1 vssd1
+ vccd1 vccd1 _02579_ sky130_fd_sc_hd__or2_1
XANTENNA__06587__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _01078_ net161 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__nand2_1
X_09627_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\] _04694_ vssd1
+ vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06839_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] _02498_ _02509_
+ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__o21ai_2
XANTENNA__06353__B1 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09558_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ net781 net241 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08509_ _03969_ _03970_ _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09489_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ net268 _04619_ net290 net222 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08307__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10402_ clknet_leaf_17_wb_clk_i net706 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08948__A3 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10333_ clknet_leaf_26_wb_clk_i net726 net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10264_ clknet_leaf_7_wb_clk_i _00256_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10195_ clknet_leaf_83_wb_clk_i _00199_ net301 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05953__X _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout380 net385 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_2
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05934__A3 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06895__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10844__519 vssd1 vssd1 vccd1 vccd1 _10844__519/HI net519 sky130_fd_sc_hd__conb_1
XFILLER_0_68_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput11 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput22 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05170_ _00849_ _00877_ _00882_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07072__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07775__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08860_ _00797_ _00959_ _00960_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nor3_1
X_07811_ _01095_ net148 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08791_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] _04147_ vssd1
+ vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__or2_1
X_07742_ _03281_ _03283_ _03296_ _03276_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__o31ai_1
X_04954_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1 vssd1 vccd1
+ vccd1 _00694_ sky130_fd_sc_hd__inv_2
XANTENNA__07127__A2 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07673_ net155 _03229_ _03230_ _03228_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09412_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _02965_ _04556_ _02963_
+ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__o22a_2
XFILLER_0_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06624_ _02285_ _02294_ _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09343_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__or2_1
X_06555_ net155 _01644_ net200 _01663_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout241_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05506_ _01207_ _01217_ _01218_ net418 net420 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__o32a_1
X_09274_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ net1 _04263_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07669__C _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06486_ _02092_ _02155_ _02153_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08225_ net5 _03703_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__and2b_1
X_05437_ _01130_ _01148_ _01149_ _01136_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__or4b_1
XFILLER_0_133_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10899__564 vssd1 vssd1 vccd1 vccd1 _10899__564/HI net564 sky130_fd_sc_hd__conb_1
X_08156_ net469 net471 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nor2_2
X_05368_ _01080_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07063__A1 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ net81 _02759_ _02760_ net98 _01635_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__o221a_4
X_08087_ _03596_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ net229 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05299_ _01009_ _01011_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07038_ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__and3_1
XANTENNA__06574__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05933__B _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ net591 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_98_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06877__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10882_ net557 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10947__587 vssd1 vssd1 vccd1 vccd1 _10947__587/HI net587 sky130_fd_sc_hd__conb_1
XFILLER_0_94_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05852__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07054__A1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10694__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05396__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10316_ clknet_leaf_41_wb_clk_i net743 net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10623__RESET_B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10247_ clknet_leaf_74_wb_clk_i _00239_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06004__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__A_N _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ clknet_leaf_23_wb_clk_i _00188_ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_117_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06580__A3 _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06332__A3 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06340_ _01723_ _02012_ _02013_ net414 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06271_ net180 _01929_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05222_ _00933_ _00934_ _00932_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__a21oi_1
X_08010_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06690__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05153_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__and2b_1
XANTENNA__07045__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07596__A2 _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05084_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\] _00808_
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\] vssd1
+ vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__and4bb_1
X_09961_ clknet_leaf_73_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[38\]
+ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08912_ net259 _04221_ vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__and2_1
X_09892_ net1112 net151 net149 _04882_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__a22o_1
X_08843_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] _04143_
+ net909 vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_51_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06020__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08774_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] net687 net238 vssd1
+ vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
X_05986_ net132 net128 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nand2_8
XFILLER_0_58_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ _03273_ _03274_ _03275_ _03278_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04937_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] vssd1
+ vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XANTENNA__08848__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06859__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ net143 _01689_ _01730_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__or3_1
XANTENNA__06859__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866__541 vssd1 vssd1 vccd1 vccd1 _10866__541/HI net541 sky130_fd_sc_hd__conb_1
XANTENNA__06865__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_06607_ _02266_ _02274_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__and3b_1
XFILLER_0_137_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07587_ net184 _01651_ net141 _01671_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a31o_1
X_09326_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ _04502_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__nand3_1
XFILLER_0_63_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06538_ net285 _01620_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__or2_2
XFILLER_0_69_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09257_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ _04454_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06469_ _02068_ _02101_ _02105_ _02107_ _02130_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08208_ _01261_ _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nand2_1
X_09188_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ _04404_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08139_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\] _03623_
+ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_116_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05928__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10101_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.buttonDetect
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.buttonPixel sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05944__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _00052_ _00643_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__06011__A2 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934_ net583 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07511__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10865_ net540 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10796_ clknet_leaf_70_wb_clk_i _00617_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06015__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06002__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05840_ _00714_ _01530_ _01533_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a21oi_2
X_05771_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\] _01469_
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__and4bb_1
X_07510_ _03066_ _03067_ _03068_ _03065_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__o31a_1
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ _03633_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07441_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] _03018_
+ _02984_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07372_ _02974_ _02975_ _02976_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06972__X _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__B1_N _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09111_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06323_ _01972_ _01991_ _01994_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09042_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04291_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a31o_1
XANTENNA__06474__C1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06254_ net456 net212 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05205_ _00916_ _00917_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] vssd1 vssd1 vccd1
+ vccd1 net1069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__dlygate4sd3_1
X_06185_ _01856_ _01865_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout204_A _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\] vssd1 vssd1 vccd1
+ vccd1 net1091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold433 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\] vssd1 vssd1
+ vccd1 vccd1 net1102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__dlygate4sd3_1
X_05136_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__nor2_1
Xhold455 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\] vssd1 vssd1
+ vccd1 vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06777__B1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold477 team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\] vssd1 vssd1 vccd1
+ vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ net461 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
X_05067_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back _00795_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select vssd1
+ vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__nor4b_4
XFILLER_0_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold488 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ net153 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout194_X net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08826_ net1126 _04141_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07741__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
X_05969_ net251 _01658_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__nand2_4
X_07708_ _01675_ _03261_ _03262_ _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06595__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ _04073_ _04107_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a41o_1
XFILLER_0_138_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07639_ _01655_ _01728_ _01874_ _03196_ net254 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05930__C _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10650_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_rs_enable
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.sck_rs_enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ clknet_leaf_60_wb_clk_i _00012_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08034__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05945__Y _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07592__C _03149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05991__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ clknet_leaf_31_wb_clk_i net879 net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10364__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06001__C _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10962__602 vssd1 vssd1 vccd1 vccd1 _10962__602/HI net602 sky130_fd_sc_hd__conb_1
X_10917_ net661 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10848_ net523 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10779_ clknet_leaf_64_wb_clk_i _00600_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07486__D _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__C1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07990_ _03532_ _03537_ _03538_ _03544_ _03531_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__o221a_1
Xfanout209 _04325_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06941_ net427 _02500_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05982__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06399__B _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09660_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\]
+ _04717_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__and3_1
X_06872_ net430 _02528_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__nor2_1
X_08611_ _04041_ _04040_ _04037_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05823_ _01513_ _01516_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__and2_1
X_09591_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ _03996_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__nand2_1
X_05754_ _01448_ _01451_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\] _03944_
+ _03713_ net463 vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__o211a_1
X_05685_ net437 net436 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout154_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07424_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] _03008_
+ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07239__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout321_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06306_ _01974_ _01976_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__or3b_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07286_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09025_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04280_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06462__A2 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__D team_07_WB.instance_to_wrap.team_07.recHEART.heartDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06237_ _01838_ _01869_ _01875_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__and4b_1
XFILLER_0_5_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold230 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] vssd1 vssd1
+ vccd1 vccd1 net899 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ net286 _01679_ _01689_ _01848_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a31o_1
Xhold241 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold263 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] vssd1 vssd1
+ vccd1 vccd1 net943 sky130_fd_sc_hd__dlygate4sd3_1
X_05119_ net299 _00830_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__nor2_1
XANTENNA__07693__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[4\]
+ vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
X_06099_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\]
+ _01781_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__or3_1
Xhold296 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\] vssd1 vssd1 vccd1
+ vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09927_ _01785_ net149 _04903_ net836 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__a22o_1
XANTENNA__10387__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ net1119 _04824_ _04860_ _04805_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08911__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ net983 _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__nand2_1
X_09789_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\] _04808_ _04812_
+ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__a21o_1
XANTENNA__05941__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10702_ clknet_leaf_66_wb_clk_i _00533_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08744__S net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06150__A1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10467__RESET_B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10633_ clknet_leaf_38_wb_clk_i _00497_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10564_ clknet_leaf_6_wb_clk_i _00432_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07650__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10495_ clknet_leaf_14_wb_clk_i _00363_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07108__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07469__A1 _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05470_ _01061_ _01096_ _01064_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06141__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06692__A2 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10137__RESET_B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ _02791_ _02792_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07071_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\] net299 _00943_ _02724_
+ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06022_ net143 _01667_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__nand2_2
XANTENNA__07794__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06601__C1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ _03525_ _03527_ _03526_ _03367_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__or4b_1
X_09712_ _04754_ _04755_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\]
+ _04730_ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a2bb2o_1
X_06924_ net174 _02511_ _02594_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07018__B _00828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07157__B1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__nand4b_1
X_06855_ _02525_ _02503_ _02497_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout271_A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05806_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] _01496_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] vssd1 vssd1
+ vccd1 vccd1 _01500_ sky130_fd_sc_hd__and3b_1
XFILLER_0_117_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09574_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] _01418_
+ _04661_ net482 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__o31a_1
XANTENNA__06380__A1 _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06786_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ _02413_ _00673_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07034__A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ net1008 _03978_ _03986_ vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_26_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05737_ _01437_ _01440_ _01439_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ _03709_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_137_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06132__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05668_ _00678_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] vssd1 vssd1 vccd1
+ vccd1 _01381_ sky130_fd_sc_hd__nor3_2
XFILLER_0_136_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07407_ _02998_ net230 _02997_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07880__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ _03753_ _03862_ net129 vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06592__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05599_ _01305_ _01306_ _01311_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07338_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\] team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07269_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ _02904_ _02907_ _01315_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[17\]
+ sky130_fd_sc_hd__a211o_1
X_09008_ net247 _04272_ _04273_ net404 net1137 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__a32o_1
XANTENNA__05001__B _00735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ clknet_leaf_80_wb_clk_i _00272_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05936__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05946__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07148__B1 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05952__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__X _02074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06123__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08327__X _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10616_ clknet_leaf_40_wb_clk_i _00480_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10547_ clknet_leaf_11_wb_clk_i _00415_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07623__A1 _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06007__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10478_ clknet_leaf_28_wb_clk_i _00346_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09318__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07926__A2 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04970_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1 vssd1 vccd1
+ vccd1 _00709_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06640_ _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06571_ _02129_ _02242_ _02243_ _02244_ _02241_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08310_ _01306_ _03682_ _03786_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05522_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _01232_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__nor2_1
X_09290_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06114__A1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ team_07_WB.instance_to_wrap.team_07.circlePixel net486 vssd1 vssd1 vccd1
+ vccd1 _03720_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_28_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06665__A2 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05453_ _01057_ _01075_ _01111_ _01160_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_131_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07862__B2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08172_ _03628_ _03648_ _03651_ _03649_ net463 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05384_ net191 _01005_ _01021_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_132_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07123_ _02764_ _02767_ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__a21o_1
XANTENNA__07614__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06417__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901__566 vssd1 vssd1 vccd1 vccd1 _10901__566/HI net566 sky130_fd_sc_hd__conb_1
XFILLER_0_3_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout117_A _01608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ net271 net269 _01638_ _02335_ _02708_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__o311a_1
XANTENNA__08413__A _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06005_ net157 net147 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_28_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07956_ _01057_ _01741_ _03371_ _03510_ net252 vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__o221a_1
X_06907_ net428 net182 _02505_ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a211o_1
X_07887_ _01078_ net158 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__or2_1
XANTENNA__08878__B1 _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06587__B _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ net1096 _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__nor2_1
X_06838_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__nand2_2
XANTENNA__06353__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ net1178 net241 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
X_06769_ _02417_ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__nor2_1
X_08508_ _03969_ _03970_ _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__and4_1
XANTENNA__07699__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09488_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04616_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_121_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05836__B1_N _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08439_ net460 _03912_ _03681_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10401_ clknet_leaf_17_wb_clk_i net682 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07605__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ clknet_leaf_25_wb_clk_i net704 net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ clknet_leaf_7_wb_clk_i _00255_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ clknet_leaf_81_wb_clk_i _00198_ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout370 net385 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_2
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_4
Xfanout392 _03024_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06344__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883__558 vssd1 vssd1 vccd1 vccd1 _10883__558/HI net558 sky130_fd_sc_hd__conb_1
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05855__B1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput12 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput23 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07057__C1 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10185__D net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ _01094_ net144 vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08790_ _04147_ _04148_ net192 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__a21oi_1
X_10818__493 vssd1 vssd1 vccd1 vccd1 _10818__493/HI net493 sky130_fd_sc_hd__conb_1
XANTENNA__06583__A1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05592__A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _01064_ net115 _03291_ _00750_ _03290_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__o221a_1
XANTENNA__06040__X _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04953_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07672_ _01680_ _02055_ _02081_ _01646_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__a22o_1
XANTENNA__06335__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ net873 _04566_ _04565_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06623_ _02280_ _02292_ _02269_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nand2_1
X_06554_ _02139_ net85 _02214_ _02149_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05505_ _01199_ _01216_ _01210_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__o21ai_1
X_09273_ net3 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ _04469_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__mux2_1
X_06485_ _01636_ _02157_ _02158_ _02109_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ net6 net1 vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__nor2_1
X_05436_ net431 _01072_ _01131_ net296 _01146_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08155_ net468 net470 vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout401_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05367_ net189 _01025_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__nor2_1
X_07106_ _01630_ _01636_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08086_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ _00814_ net476 vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__o21a_1
XANTENNA__07063__A2 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05298_ net189 _01004_ _01010_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07037_ _02677_ _02681_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__or2_2
XFILLER_0_12_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06023__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06598__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ _04257_ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07939_ _01078_ net198 net187 _01084_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_3_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ net590 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_3_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06326__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__B1 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05007__A _00738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] _04682_ vssd1
+ vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__or2_1
X_10881_ net556 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_39_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07222__A _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08752__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07054__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10315_ clknet_leaf_41_wb_clk_i net736 net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08075__A_N net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10246_ clknet_leaf_71_wb_clk_i _00238_ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10177_ clknet_leaf_24_wb_clk_i _00187_ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07109__A3 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07132__A _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06270_ net138 _01926_ _01928_ net156 _01946_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05221_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00934_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05152_ _00861_ _00864_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05083_ _00705_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\] vssd1
+ vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__or3_1
X_09960_ clknet_leaf_82_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[29\]
+ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08911_ net435 _01400_ _01403_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__a31o_1
X_09891_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] _01775_ vssd1
+ vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__xnor2_1
X_08842_ net964 _04143_ _04181_ vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_51_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__A _02930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] net702 net237 vssd1
+ vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__mux2_1
XANTENNA__06020__A3 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05985_ net133 net121 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__nor2_4
XFILLER_0_109_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout184_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ _03273_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04936_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] vssd1 vssd1
+ vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07505__B1 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _02734_ _03181_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout351_A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout449_A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ net134 net125 _01936_ _02275_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__or4_1
XFILLER_0_88_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07586_ net256 net179 _02151_ _01663_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o31a_1
XFILLER_0_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09325_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04499_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a31o_1
XANTENNA__07042__A _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06537_ _02208_ _02210_ _02207_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout237_X net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10907__572 vssd1 vssd1 vccd1 vccd1 _10907__572/HI net572 sky130_fd_sc_hd__conb_1
X_09256_ net227 _04456_ _04457_ net405 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06468_ _02119_ _02126_ _02133_ _01625_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06881__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08207_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] _03682_
+ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05419_ _01034_ _01036_ _01039_ _01099_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_43_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09187_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ _04404_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__or2_1
XANTENNA__07696__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06399_ net176 _01732_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__nand2_4
XFILLER_0_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ _03624_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__A3 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08069_ net454 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__and2b_1
X_10100_ clknet_3_4_0_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.stageDetect
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.stagePixel
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout97_A _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _00051_ _00047_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05944__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08747__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10933_ net582 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07511__A3 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net539 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_39_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10795_ clknet_leaf_70_wb_clk_i _00616_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05959__X _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07887__A _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07680__C1 _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06015__B net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10229_ clknet_leaf_79_wb_clk_i _00233_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06031__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05770_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] vssd1 vssd1 vccd1
+ vccd1 _01469_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07499__C1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] _03018_
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06710__A1 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05513__A2 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07371_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02969_
+ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04347_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__and2_1
X_06322_ _01972_ _01983_ _01994_ _01997_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09041_ net247 _04296_ _04297_ net407 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__a32o_1
XANTENNA__06474__B1 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06253_ net212 _01926_ _01929_ net194 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05204_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00917_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold401 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06184_ net175 net120 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10364__SET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold412 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\] vssd1 vssd1
+ vccd1 vccd1 net1081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] vssd1 vssd1
+ vccd1 vccd1 net1092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] vssd1 vssd1
+ vccd1 vccd1 net1103 sky130_fd_sc_hd__dlygate4sd3_1
X_05135_ _00845_ _00847_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold445 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold456 team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\] vssd1 vssd1 vccd1
+ vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] vssd1 vssd1
+ vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold478 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ net461 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
X_05066_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _00793_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__or2_2
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_A _00807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ net998 net153 _04871_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a21o_1
XANTENNA__06529__A1 _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07037__A _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _04141_
+ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06544__A4 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ net1130 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__mux2_1
X_05968_ _01489_ net215 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__nand2_2
X_04919_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
X_07707_ _02040_ _02877_ _01744_ _01795_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a211o_1
X_05899_ _01591_ _01592_ _01574_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a21boi_4
X_08687_ _04046_ _04109_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07638_ _01644_ _01675_ _01742_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_68_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07569_ _01611_ _02332_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09308_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ _04491_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and2_1
XANTENNA__05004__B net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10580_ clknet_leaf_60_wb_clk_i _00011_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07500__A _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ net227 _04443_ _04445_ net406 net786 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05020__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06768__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05955__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05991__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ clknet_leaf_31_wb_clk_i _00093_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08390__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05961__Y _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05690__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10916_ net660 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08693__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08209__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10847_ net522 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_39_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10778_ clknet_leaf_65_wb_clk_i _00599_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06456__B1 _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08225__B _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06671__D _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06026__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06940_ _02522_ _02596_ _02605_ _02610_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06032__Y _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05982__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06871_ _02533_ _02541_ net134 _02526_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05822_ _01492_ _01493_ _01501_ _01515_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__o31a_4
XFILLER_0_59_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08610_ _00689_ _01201_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__xnor2_1
X_09590_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] vssd1 vssd1 vccd1 vccd1
+ _04671_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06931__B2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05753_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] vssd1 vssd1 vccd1
+ vccd1 _01452_ sky130_fd_sc_hd__or3_1
X_08541_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08472_ _03770_ _03942_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__and3_1
X_05684_ net437 net436 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07423_ _03008_ net477 _03007_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[14\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07354_ _02961_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_98_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07239__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06305_ _01978_ _01979_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__and3b_1
XANTENNA__07320__A _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07285_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ _02914_ _02917_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[11\]
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_135_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout314_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ _04283_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06236_ net100 _01671_ _01874_ _01914_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10454__Q team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net127
+ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__xnor2_1
Xhold231 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout102_X net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__dlygate4sd3_1
X_05118_ net447 team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] _00685_ vssd1
+ vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__and3b_1
XFILLER_0_40_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold275 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[1\] vssd1
+ vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__dlygate4sd3_1
X_06098_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] _01780_
+ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold286 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] _01784_
+ net152 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__or3_1
X_05049_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00780_ vssd1 vssd1
+ vccd1 vccd1 _00781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09857_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] _04858_ vssd1
+ vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08808_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] _04154_ vssd1 vssd1
+ vccd1 vccd1 _04160_ sky130_fd_sc_hd__or4_4
X_10985__625 vssd1 vssd1 vccd1 vccd1 _10985__625/HI net625 sky130_fd_sc_hd__conb_1
X_09788_ _01768_ _04810_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__and3_1
X_08739_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ net233 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10701_ clknet_leaf_66_wb_clk_i _00532_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06150__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10632_ clknet_leaf_40_wb_clk_i _00496_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10563_ clknet_leaf_8_wb_clk_i _00431_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05021__Y _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10494_ clknet_leaf_16_wb_clk_i _00362_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07650__A2 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06677__B1 _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06429__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07070_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\]
+ net446 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05298__C _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06021_ net138 _01708_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05404__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07972_ _01113_ net172 net252 vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__o21ai_1
X_09711_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] _04752_ _04731_
+ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__o21ai_1
X_06923_ net186 _02508_ _02577_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a21oi_1
X_10969__609 vssd1 vssd1 vccd1 vccd1 _10969__609/HI net609 sky130_fd_sc_hd__conb_1
XANTENNA__07157__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09642_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__or4_1
X_06854_ _02499_ _02504_ _02524_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a21bo_1
X_05805_ _01495_ _01496_ _01498_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_96_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06785_ _02410_ _02414_ net93 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a21oi_1
X_09573_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04629_ _04657_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__or3_2
XFILLER_0_117_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08524_ _03985_ _03976_ _03984_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__or3b_1
X_05736_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ _00652_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06668__B1 _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08455_ net486 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ net488 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] vssd1 vssd1
+ vccd1 vccd1 _03928_ sky130_fd_sc_hd__or4b_1
X_05667_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] vssd1 vssd1 vccd1
+ vccd1 _01380_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_93_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__04945__Y _00685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06132__A2 _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07406_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\]
+ _02994_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08386_ net462 _03859_ _03861_ _03749_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_82_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05598_ _01303_ _01304_ _01302_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07337_ _02947_ _02949_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ _01315_ _02907_ _02908_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[16\]
+ sky130_fd_sc_hd__nor3_1
X_09007_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06219_ net97 _01878_ _01885_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05776__Y _01475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ _01739_ _02036_ _02836_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07991__Y team_07_WB.instance_to_wrap.team_07.recGen.circleDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05946__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] _01779_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] vssd1 vssd1 vccd1
+ vccd1 _04893_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_109_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05952__B _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08755__S net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06674__A3 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05399__B _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10615_ clknet_leaf_40_wb_clk_i _00479_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10546_ clknet_leaf_11_wb_clk_i _00414_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07623__A2 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10477_ clknet_leaf_28_wb_clk_i _00345_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06304__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09128__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06570_ _02050_ _02114_ _02134_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06974__A _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05521_ _01219_ _01232_ _01233_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07789__B _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06114__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06693__B _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ team_07_WB.instance_to_wrap.team_07.circlePixel net486 vssd1 vssd1 vccd1
+ vccd1 _03719_ sky130_fd_sc_hd__and2b_1
X_05452_ _01163_ _01164_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ net53 _03628_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05383_ _01001_ net189 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_132_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07122_ _02768_ _02773_ _02775_ _02277_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06417__A3 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06283__D1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07053_ net86 net249 _01639_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06004_ net156 net147 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ net158 _03375_ _03458_ _03462_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__o31a_1
XANTENNA__08327__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ net428 net182 _02517_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__o21ai_1
X_07886_ _01078_ net158 vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__nor2_1
X_09625_ _04664_ _04693_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06837_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__and2_1
XANTENNA__07550__A1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06353__A2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09556_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ net773 net241 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
X_06768_ net426 net271 _02413_ _02439_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08507_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__and4bb_1
X_05719_ net479 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ _00822_ _01429_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09487_ net921 net204 _04618_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__o21a_1
X_06699_ net253 _02014_ _02048_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08438_ _00730_ _01284_ _03689_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10099__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08369_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] _03842_ _03843_
+ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ clknet_leaf_17_wb_clk_i net708 net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_132_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07605__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05616__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ clknet_leaf_25_wb_clk_i net703 net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05439__S _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ clknet_leaf_7_wb_clk_i _00254_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06124__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ clknet_leaf_82_wb_clk_i _00197_ net301 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05963__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06411__X _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout360 net385 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_2
Xfanout371 net373 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout382 net384 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_4
Xfanout393 _00968_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_4
XANTENNA__08869__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06130__Y _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06344__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
Xinput35 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10529_ clknet_leaf_31_wb_clk_i _00397_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06034__A _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07740_ net263 _03285_ _03294_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__or3_1
XANTENNA__05592__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04952_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
X_07671_ net107 net165 net162 _01678_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a22o_1
XANTENNA__06335__A2 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _04556_ vssd1 vssd1 vccd1
+ vccd1 _04566_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06622_ _01714_ _01742_ _02294_ _02293_ _02267_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09341_ net223 _04515_ _04516_ net399 net863 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a32o_1
X_06553_ _02085_ _02131_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05504_ _01203_ _01211_ _01212_ _01214_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a31o_1
X_09272_ _04420_ _04422_ _04466_ _04468_ _04421_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a2111o_1
X_06484_ _02057_ _02155_ _02153_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ _03700_ _03701_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__o21ai_2
X_05435_ _01141_ _01142_ _01143_ _01147_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__or4b_1
XANTENNA__07048__B1 _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ net468 net470 vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__and2_1
X_05366_ _00990_ _01074_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__or2_2
XFILLER_0_114_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07105_ _01636_ _02197_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__nor2_1
XANTENNA__06952__C_N team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08085_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ net229 _03595_ net897 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__a22o_1
XANTENNA__07063__A3 _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05297_ net426 _00998_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07036_ _02111_ _02687_ _02690_ _02685_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_77_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08987_ _04250_ _04251_ _04254_ _04256_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _01692_ _03492_ _03490_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_3_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07869_ net277 net393 _01063_ _03350_ _03423_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_123_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _00697_ _04680_ _04682_ _04665_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a22oi_1
X_10880_ net555 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09539_ _04650_ net910 net220 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05958__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11019__642 vssd1 vssd1 vccd1 vccd1 _11019__642/HI net642 sky130_fd_sc_hd__conb_1
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10314_ clknet_leaf_41_wb_clk_i net740 net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05964__Y _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ clknet_leaf_71_wb_clk_i _00237_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07892__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07211__B1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ clknet_leaf_23_wb_clk_i _00186_ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10850__525 vssd1 vssd1 vccd1 vccd1 _10850__525/HI net525 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
XFILLER_0_135_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07514__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload5_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07132__B _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08475__C1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06971__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05220_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00933_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05868__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06690__C net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05151_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07045__A3 _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06253__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05082_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__and3_1
XANTENNA__06253__B2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08910_ net259 _04220_ vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ net850 net151 net149 _04881_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a22o_1
XANTENNA__05835__B1_N _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] _01457_
+ _04143_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__or3_1
X_08772_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\] net783 net239 vssd1
+ vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
X_05984_ net159 net147 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__or2_4
X_07723_ _01597_ _01604_ _01105_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__a21oi_1
X_04935_ net426 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout177_A _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _01730_ _02765_ _03160_ _03211_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_95_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10373__RESET_B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06605_ net107 _01935_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07585_ _02107_ _02164_ net87 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout344_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09324_ net225 _04504_ _04505_ net401 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a32o_1
XANTENNA__05114__Y _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06536_ _02178_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ _04454_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06467_ _02060_ _02092_ _02090_ _02068_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ _03683_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05778__A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05418_ _01017_ _01033_ _01041_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__or3_1
X_09186_ net207 _04403_ _04405_ net403 net1044 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a32o_1
X_06398_ _02071_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__inv_2
XANTENNA__08769__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05349_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] net431 vssd1
+ vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__nor2_2
X_08137_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ net392 net295 net1181 _03587_ vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07019_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\]
+ net447 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
X_10834__509 vssd1 vssd1 vccd1 vccd1 _10834__509/HI net509 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_8_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ _00050_ _00046_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10953__593 vssd1 vssd1 vccd1 vccd1 _10953__593/HI net593 sky130_fd_sc_hd__conb_1
XANTENNA__07744__A1 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10932_ net581 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_86_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06294__A1_N net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10863_ net538 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_13_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08763__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10794_ clknet_leaf_70_wb_clk_i _00615_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07520__X _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07887__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07680__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07983__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__B2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891__647 vssd1 vssd1 vccd1 vccd1 net647 _10891__647/LO sky130_fd_sc_hd__conb_1
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05994__B1 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10228_ clknet_leaf_73_wb_clk_i _00232_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06312__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10159_ clknet_leaf_18_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold2 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06031__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07499__B1 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06710__A2 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02969_
+ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06321_ _01981_ _01996_ _01995_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09040_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06252_ _01926_ _01927_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__nand2_2
XFILLER_0_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05203_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00916_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06183_ net174 net120 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_96_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold402 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] vssd1 vssd1
+ vccd1 vccd1 net1071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] vssd1 vssd1
+ vccd1 vccd1 net1082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05134_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold424 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] vssd1 vssd1
+ vccd1 vccd1 net1093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] vssd1 vssd1
+ vccd1 vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ net461 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
X_05065_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up vssd1 vssd1
+ vccd1 vccd1 _00794_ sky130_fd_sc_hd__or2_1
Xhold479 team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] _04870_ vssd1
+ vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_70_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06529__A2 _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _04141_ _04170_ net193 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07037__B _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08755_ net1174 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ net233 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout461_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05967_ net256 net212 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
X_07706_ _01735_ _01901_ net184 vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__o21a_1
X_04918_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
X_08686_ net455 _04105_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a21oi_1
X_05898_ _01565_ _01569_ _01570_ _01573_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07637_ _03152_ _03178_ _03194_ _03099_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_68_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07568_ _02150_ _02191_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09307_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ _04491_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__or2_1
X_06519_ _02153_ _02189_ _02190_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_75_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07499_ net94 _02348_ _02343_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09238_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__inv_2
XANTENNA__07500__B _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05301__A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04391_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06116__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05020__B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08612__A _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06768__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05955__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07178__C1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07717__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ clknet_leaf_33_wb_clk_i _00092_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08758__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05971__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10224__RESET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05690__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10915_ net659 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
X_10846_ net521 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__05900__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10777_ clknet_leaf_65_wb_clk_i _00598_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07545__A1_N _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05211__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07956__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856__531 vssd1 vssd1 vccd1 vccd1 _10856__531/HI net531 sky130_fd_sc_hd__conb_1
XANTENNA__05865__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06042__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07708__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05982__A3 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ _02535_ _02540_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05821_ _01494_ _01497_ _01514_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07144__Y _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ _03628_ _03650_ net145 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09072__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05752_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] _01450_ vssd1 vssd1
+ vccd1 vccd1 _01451_ sky130_fd_sc_hd__or4b_1
X_08471_ net484 net487 _03710_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__or3b_1
X_05683_ net437 net436 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07422_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ _03004_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07601__A _03070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07353_ _00708_ _00816_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06304_ net198 _01977_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__B _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07284_ _02917_ _02918_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[10\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_135_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09023_ net247 _04282_ _04284_ net404 net947 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__a32o_1
X_06235_ net91 _01670_ _01706_ _01912_ _01913_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__o32a_1
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 _00094_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__dlygate4sd3_1
X_06166_ _01832_ _01836_ _01838_ _01846_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_113_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__dlygate4sd3_1
X_05117_ _00685_ _00828_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__and2_1
Xhold265 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[22\]
+ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__dlygate4sd3_1
X_06097_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\]
+ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__or3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold276 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06223__Y _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold287 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__RESET_B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09925_ net976 _01784_ _04870_ _04902_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__o31ai_1
X_05048_ _00768_ _00769_ _00770_ _00779_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__a31o_1
Xhold298 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\] vssd1 vssd1
+ vccd1 vccd1 net967 sky130_fd_sc_hd__dlygate4sd3_1
X_09856_ _04827_ _04859_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__nor2_1
X_08807_ net193 _04159_ vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__nor2_1
XANTENNA__06383__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09787_ _00657_ _04803_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__nor2_2
X_06999_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _02654_
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ net1133 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__mux2_1
XANTENNA__07537__D_N _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08669_ _04080_ _04095_ _04084_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o21ai_1
X_10700_ clknet_leaf_66_wb_clk_i _00531_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05015__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05894__C1 _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ clknet_leaf_39_wb_clk_i _00495_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07635__B1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10562_ clknet_leaf_9_wb_clk_i _00430_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06127__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10493_ clknet_leaf_16_wb_clk_i _00361_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05966__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06414__X _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06374__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06126__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06677__A1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10927__576 vssd1 vssd1 vccd1 vccd1 _10927__576/HI net576 sky130_fd_sc_hd__conb_1
X_10829_ net504 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_138_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06429__A1 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10897__653 vssd1 vssd1 vccd1 vccd1 net653 _10897__653/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_93_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06020_ net106 net141 net167 net201 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a31o_2
XFILLER_0_112_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07929__A1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07929__B2 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06601__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ _03377_ _03405_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10146__RESET_B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] _04752_ vssd1
+ vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__and2_1
X_06922_ _02591_ _02592_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__or2_1
XANTENNA__07157__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__or4b_1
XFILLER_0_93_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05168__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06853_ _02499_ _02504_ _02507_ net186 _02523_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05804_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] _01486_
+ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__nand2_1
X_09572_ net482 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04657_ _04660_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a31o_1
X_06784_ _02431_ _02454_ _02455_ _02428_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05116__A _00685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ _03983_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05735_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\] _00787_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_65_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout257_A _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06668__B2 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ _03667_ _03826_ _03923_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04955__A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05666_ net415 _00676_ _00677_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_137_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07405_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] _02994_
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] vssd1 vssd1 vccd1
+ vccd1 _02997_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_102_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08385_ _03718_ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_82_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05597_ _01302_ _01303_ _01304_ _01309_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_82_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07336_ _02414_ _02948_ _01175_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09006_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06218_ _01894_ _01895_ _01897_ _01889_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07198_ _02773_ _02846_ _02781_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06149_ net103 _01828_ net210 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05946__A3 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ net1106 net152 net150 _04892_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a22o_1
XANTENNA__07148__A2 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ net243 _04845_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10614_ clknet_leaf_40_wb_clk_i _00478_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07608__B1 _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07084__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10545_ clknet_leaf_10_wb_clk_i _00413_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05967__Y _01661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10476_ clknet_leaf_28_wb_clk_i _00344_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06347__B1 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06898__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05520_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01219_ _01232_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07789__C _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05451_ _01042_ _01068_ _01102_ _01020_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__o22a_1
XANTENNA__05322__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08170_ net463 _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05382_ _00970_ _01063_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__nand2_2
XFILLER_0_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07075__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _01635_ _02757_ _02769_ _02774_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10398__RESET_B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06283__C1 _01959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07052_ _02677_ _02691_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06003_ net216 net195 _01682_ _01695_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__o31a_2
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07954_ _01057_ _01658_ _03369_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__a21o_1
XANTENNA__08327__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ net428 net182 net171 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__o2bb2a_1
X_07885_ net262 _03285_ _03413_ _03439_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout374_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _04666_ _04692_ _04693_ _04664_ net1048 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a32o_1
X_06836_ net427 _02506_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__nor2_1
XANTENNA__07550__A2 _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ net217 _04605_ net881 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_06767_ net275 net425 net273 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_104_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08506_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__and3_1
X_05718_ net476 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09486_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ net268 _04617_ net290 net222 vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a221o_1
X_06698_ net174 _02274_ net253 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05133__X _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08437_ _00711_ _00727_ _03717_ _03910_ _00048_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05649_ _01360_ _01361_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07996__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08368_ _00729_ _01380_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__nand2_1
XANTENNA__09055__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07319_ _01190_ _01192_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08263__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08299_ net5 _00663_ _03703_ _03705_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a41o_1
XFILLER_0_116_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10330_ clknet_leaf_24_wb_clk_i net685 net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_108_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10261_ clknet_leaf_7_wb_clk_i _00253_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10192_ clknet_leaf_81_wb_clk_i net1095 net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05963__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_128_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07236__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_4
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06329__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08869__A2 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout394 _00943_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_2
XFILLER_0_69_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__B1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06501__B1 _02149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05978__X _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05203__B _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05855__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07057__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10528_ clknet_leaf_31_wb_clk_i _00396_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06804__B2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ clknet_leaf_27_wb_clk_i net1050 net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06034__B _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07146__A _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06050__A _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04951_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
X_07670_ net104 _02277_ _03173_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o21a_1
X_06621_ _01698_ _02021_ net255 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09340_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a31o_1
X_06552_ _01618_ net249 _02196_ net261 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05503_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ _01215_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__xnor2_1
X_09271_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ _04467_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__or3b_1
XFILLER_0_59_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06483_ _02155_ _02156_ _02153_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel _00728_ team_07_WB.instance_to_wrap.team_07.buttonPixel
+ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05434_ _00982_ _01027_ _01091_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08153_ net468 _00717_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__and2_1
X_05365_ net393 _01056_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__nand2_4
XFILLER_0_16_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout122_A _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07104_ net81 _02756_ _02757_ _01635_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__o211a_4
XFILLER_0_70_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[6\]
+ net229 _03595_ net878 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06225__A _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05296_ _01001_ _01008_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07035_ _02688_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_77_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06023__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__or4_1
X_07937_ _03487_ _03491_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07868_ _00968_ _01058_ _02106_ _00749_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_3_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__A2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09607_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\]
+ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and3_1
X_06819_ net113 _02477_ _02478_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07799_ _03340_ _03346_ _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__or3_2
X_09538_ net289 _04645_ _04649_ net267 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05638__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09469_ net900 net202 _04607_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05023__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10249__RESET_B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07039__A1 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05958__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06406__Y _02080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ clknet_leaf_41_wb_clk_i net746 net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05974__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05470__B1 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ clknet_leaf_71_wb_clk_i _00236_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07211__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ clknet_leaf_22_wb_clk_i _00185_ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06905__A2_N net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
Xfanout191 _00990_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05980__Y team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07514__A2 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05525__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05150_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] _00862_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_4
XFILLER_0_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05081_ _00807_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ sky130_fd_sc_hd__inv_2
XFILLER_0_110_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05461__B1 _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08840_ _04143_ _04180_ _04144_ vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06051__Y _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08950__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] net733 net239 vssd1
+ vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05983_ net158 net146 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__nor2_4
XFILLER_0_58_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06961__B1 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _01064_ net115 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__nor2_1
X_04934_ net425 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07604__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _03063_ _03064_ _03210_ _03209_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__o31a_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_X clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06604_ _01651_ _01936_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__nor2_4
XFILLER_0_76_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07584_ _02232_ _03142_ _02830_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__o21ba_1
X_09323_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ _04502_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__nand2_1
X_06535_ net263 net271 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__or2_2
XANTENNA__07269__A1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout337_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ _04454_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or2_1
XANTENNA__07674__D1 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06466_ _00752_ _02030_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__or2_2
XFILLER_0_91_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ net417 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _01258_
+ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05417_ _00668_ _01055_ _01129_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__a21oi_1
X_09185_ _04404_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06397_ net164 _02069_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03621_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or4_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05348_ net191 _01000_ _01004_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__or3_2
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08067_ net454 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05279_ _00979_ _00987_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07018_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] _00828_ vssd1 vssd1
+ vccd1 vccd1 _02673_ sky130_fd_sc_hd__nor2_2
XANTENNA__08170__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873__548 vssd1 vssd1 vccd1 vccd1 _10873__548/HI net548 sky130_fd_sc_hd__conb_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07744__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08969_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] net822
+ net444 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XANTENNA__05018__B net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ net580 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10862_ net537 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10793_ clknet_leaf_70_wb_clk_i _00614_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05969__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10083__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09728__X _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05443__B1 _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05994__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ clknet_leaf_79_wb_clk_i _00231_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09463__X _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05991__X _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ clknet_leaf_19_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[5\]
+ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10089_ clknet_leaf_66_wb_clk_i _00147_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07499__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06320_ net177 _01973_ _01984_ _01986_ _01976_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a41o_1
X_06251_ _01927_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__inv_2
XANTENNA__07671__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07671__B2 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06046__Y _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05202_ _00907_ _00914_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06182_ _01858_ _01860_ _01861_ _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_96_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold403 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold414 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05133_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\]
+ _00843_ _00840_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux4_2
XFILLER_0_128_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold425 team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] vssd1 vssd1 vccd1
+ vccd1 net1094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold436 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold447 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\] vssd1 vssd1
+ vccd1 vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09941_ net461 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
Xhold469 net56 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__dlygate4sd3_1
X_05064_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right vssd1
+ vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ net333 _01790_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07187__B1 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08823_ net805 _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__nand2_1
XANTENNA__06934__B1 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08754_ net1037 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
X_05966_ net256 _01659_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__nor2_4
XFILLER_0_135_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07705_ net165 net102 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__nand2_1
X_04917_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08685_ _04049_ _04073_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__and3_1
X_05897_ _01562_ net147 _01572_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07636_ _02061_ _03193_ _03165_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06162__A1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06162__B2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07567_ _02217_ _02223_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout242_X net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09306_ net226 _04490_ _04492_ net398 net1032 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06518_ _02108_ _02150_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07498_ _00943_ _02250_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__and3b_1
XFILLER_0_35_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09237_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04418_ _04435_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06449_ _01686_ _01703_ _01722_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__or3_1
XFILLER_0_111_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09168_ net207 _04390_ _04392_ net403 net800 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08119_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\] vssd1
+ vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05795__Y _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04318_ _04333_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07178__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ clknet_leaf_21_wb_clk_i _00009_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05728__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05971__B net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input15_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10914_ net658 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_10845_ net520 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10776_ clknet_leaf_65_wb_clk_i _00597_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05211__B _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__A2 _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06042__B _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05820_ _01495_ _01496_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__nor2_1
XANTENNA__07154__A _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05751_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] _01449_ vssd1 vssd1
+ vccd1 vccd1 _01450_ sky130_fd_sc_hd__nor4_1
XFILLER_0_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08470_ _00729_ _03940_ _03941_ _03738_ net484 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a311o_1
XFILLER_0_106_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05682_ _01318_ _01393_ _01394_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__nand3_1
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07421_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ _03003_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\] vssd1
+ vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07352_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\] _02958_
+ _02960_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__or4_2
XFILLER_0_9_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06303_ net213 _01967_ _01968_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__or3_1
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07283_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09022_ _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06234_ net114 _01880_ _01911_ net91 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold200 _00484_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__dlygate4sd3_1
X_06165_ _01839_ _01845_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout202_A _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__dlygate4sd3_1
X_05116_ _00685_ _00828_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__nor2_1
Xhold244 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\] vssd1 vssd1
+ vccd1 vccd1 net913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06096_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] _01778_
+ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__or2_1
Xhold266 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] vssd1 vssd1
+ vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _01784_ net152 net976 vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__o21ai_1
X_05047_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\]
+ _00777_ _00778_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06520__X _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ net243 _04858_ _04857_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input7_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net1081 _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06383__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06998_ _02655_ _02656_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__and3_1
X_09786_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nand2_1
XANTENNA__10704__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07064__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__mux2_1
X_05949_ net210 _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__nand2_1
XANTENNA__07999__A team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07332__A0 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ _04089_ _04092_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07619_ net250 _01731_ _02271_ _03114_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__a211o_1
X_08599_ _03624_ _04033_ _03626_ vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ clknet_leaf_39_wb_clk_i _00494_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09981__SET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06408__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10561_ clknet_leaf_8_wb_clk_i _00429_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07635__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922__666 vssd1 vssd1 vccd1 vccd1 net666 _10922__666/LO sky130_fd_sc_hd__conb_1
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06127__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10492_ clknet_leaf_16_wb_clk_i _00360_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10879__554 vssd1 vssd1 vccd1 vccd1 _10879__554/HI net554 sky130_fd_sc_hd__conb_1
XANTENNA__06143__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08769__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__B1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05206__B _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06677__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10828_ net503 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_89_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06429__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10759_ clknet_leaf_60_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[6\]
+ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05876__B _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07929__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06053__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06601__A2 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _01692_ _03385_ _03524_ _03523_ net106 vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_39_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05892__A _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ net427 net182 _02509_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__and3_1
X_09640_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _04702_ _00761_
+ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__o21ai_1
X_06852_ net427 net182 _02506_ _02517_ _02522_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__o311a_1
XANTENNA__05168__A2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10186__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05803_ _01495_ _01496_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ _04657_ _04625_ _04612_ _01421_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__and4b_1
X_06783_ _02426_ _02450_ _02451_ _02448_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__o2bb2a_1
X_08522_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\] _03983_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05116__B _00828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05734_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\] _01437_ _01438_
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\]
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08708__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ _03925_ _03630_ _03631_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__or3b_1
X_05665_ _01371_ _01377_ net439 _01322_ _01370_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_137_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07404_ net1001 _02994_ _02996_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_08384_ _03739_ _03805_ _03723_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05596_ _01303_ _01304_ _01307_ _01308_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_102_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07617__A1 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ _02413_ _02947_ _00965_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07266_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10100__CLK clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ _04253_ net247 _04271_ net404 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06217_ net101 _01824_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__o21bai_1
X_07197_ _02040_ _02775_ _02836_ _02848_ _02767_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07059__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10991__631 vssd1 vssd1 vccd1 vccd1 _10991__631/HI net631 sky130_fd_sc_hd__conb_1
X_06148_ net177 _01723_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__nand2_4
XFILLER_0_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06079_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] _01763_ _01764_
+ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__and4_1
X_09907_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] _01779_
+ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__xnor2_1
X_09838_ net264 _04845_ _04846_ net243 net1069 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09769_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_126_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10234__SET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05026__B _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07856__B2 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06513__D1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10613_ clknet_leaf_40_wb_clk_i _00477_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07608__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10544_ clknet_leaf_11_wb_clk_i _00412_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07084__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ clknet_leaf_27_wb_clk_i _00343_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06044__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05983__Y _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07847__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05450_ _01009_ _01076_ _01103_ _01069_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__o22a_1
XANTENNA__08962__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06048__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05381_ net296 _01062_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_132_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07120_ net88 _02109_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10975__615 vssd1 vssd1 vccd1 vccd1 _10975__615/HI net615 sky130_fd_sc_hd__conb_1
X_07051_ _01902_ _02087_ _02695_ _02705_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a31o_1
XANTENNA__06283__B1 _01957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06054__Y _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06002_ net168 net104 _01693_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__X team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06511__A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ net272 _03355_ _03356_ _03506_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06904_ _02534_ _02574_ _02532_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a21oi_1
X_07884_ _03285_ _03438_ _03282_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09623_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ _04688_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__nand3_1
X_06835_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__nor2_1
X_09554_ net881 net202 _04656_ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__o21a_1
X_06766_ net90 _02413_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_104_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07342__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__nor4_1
X_05717_ _01412_ _01413_ _01425_ _01428_ net242 vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_19_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06697_ _02214_ _02258_ _02362_ net261 _02190_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a221o_1
X_09485_ _04613_ _04616_ _00667_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08436_ _03835_ _03909_ net488 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21o_1
X_05648_ _00678_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01359_ vssd1
+ vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__a31o_1
XANTENNA__08872__S net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08367_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] _01270_ _01296_
+ _01302_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel vssd1 vssd1
+ vccd1 vccd1 _03843_ sky130_fd_sc_hd__a41o_1
XFILLER_0_135_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05579_ _01281_ _01289_ _01290_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04972__Y _00711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07318_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08298_ team_07_WB.instance_to_wrap.team_07.heartPixel _03775_ net487 vssd1 vssd1
+ vccd1 vccd1 _03776_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05077__B2 _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07249_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06405__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ clknet_leaf_7_wb_clk_i _00252_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10766__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ clknet_leaf_81_wb_clk_i _00195_ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08112__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout340 net350 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout351 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07236__B _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05308__Y _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06329__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_2
Xfanout395 net398 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_2
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07829__A1 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07829__B2 _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07057__A2 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_1
XFILLER_0_52_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput26 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput37 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10527_ clknet_leaf_30_wb_clk_i _00395_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ clknet_leaf_13_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_back
+ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06568__A1 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10389_ clknet_leaf_2_wb_clk_i net819 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_36_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06331__A team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07146__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04950_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06050__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__S _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06620_ _02280_ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__and2_1
X_06551_ _02220_ _02222_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05502_ net418 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__nand2b_1
X_09270_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04420_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__or4b_1
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06482_ net102 _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08221_ team_07_WB.instance_to_wrap.team_07.heartPixel team_07_WB.instance_to_wrap.team_07.labelPixel\[1\]
+ _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05433_ _01059_ _01060_ _01144_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11003__637 vssd1 vssd1 vccd1 vccd1 _11003__637/HI net637 sky130_fd_sc_hd__conb_1
XFILLER_0_117_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08152_ net471 _03635_ _03637_ _03634_ vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__a22o_1
X_05364_ net433 _01049_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__or2_2
XANTENNA__06506__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload54_A clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ _02249_ net81 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08083_ net878 net229 _03595_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05295_ net421 net422 _00988_ _00980_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout115_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06225__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07034_ _02085_ _02185_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06241__A _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or4b_1
XFILLER_0_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07936_ net252 _03475_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ net269 _03392_ _03395_ _03396_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__or4_1
XFILLER_0_98_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__04967__Y _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\]
+ _04675_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06818_ _02478_ _02488_ net120 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__a21o_1
XANTENNA__05007__D _00743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08168__A _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07798_ _03347_ _03350_ _03351_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09537_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _01420_
+ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__or2_1
X_06749_ _00672_ net146 net154 net423 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09468_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ net265 net287 net217 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07800__A _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08419_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] _00704_
+ _03646_ _03893_ _03630_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a41o_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09399_ _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08236__A1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06135__B _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ clknet_leaf_41_wb_clk_i net724 net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_105_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10243_ clknet_leaf_78_wb_clk_i _00235_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05974__B net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ clknet_leaf_23_wb_clk_i _00184_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_121_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06151__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout170 _01668_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
Xfanout181 _01532_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout192 net193 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
XANTENNA__06707__D1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07683__C1 _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08227__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05868__C _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05080_ team_07_WB.EN_VAL_REG _00065_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__nand2_8
XFILLER_0_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06061__A _00685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08950__A2 _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] net744 net239 vssd1
+ vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
X_05982_ net157 net130 net124 net138 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_72_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07721_ _03274_ _03275_ _03273_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__o21bai_1
X_04933_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07652_ _01904_ _02278_ _03188_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__o21a_1
XANTENNA__07604__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06713__A1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05516__A2 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06603_ _02275_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__inv_2
X_07583_ _01655_ _01717_ _01828_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09322_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ _04502_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__or2_1
X_06534_ _02129_ _02150_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09253_ net228 _04453_ _04455_ net406 net939 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06465_ _00752_ _02030_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout232_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10729__RESET_B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\]
+ _00730_ _01260_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__and4_1
X_05416_ _00966_ _01089_ _01128_ _01064_ _01075_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09184_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__and3_1
X_06396_ _01676_ _01688_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05140__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03621_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nor2_1
X_05347_ _01000_ net188 _01021_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout118_X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ net391 net293 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ _03586_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_116_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07013__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05278_ net190 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07017_ net903 _02672_ _02670_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08968_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] net791
+ net444 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
X_07919_ _03305_ _03445_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__nor2_1
X_08899_ net479 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\] vssd1
+ vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__and3_1
X_10930_ net579 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__07901__B1 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10861_ net536 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_21_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06180__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10792_ clknet_leaf_70_wb_clk_i _00613_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05969__B _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__A2 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05985__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10226_ clknet_leaf_73_wb_clk_i _00230_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05209__B _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ clknet_leaf_16_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06943__A1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_50_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07705__A net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ clknet_leaf_66_wb_clk_i _00146_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07499__A2 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_X clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06250_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] net456 vssd1 vssd1
+ vccd1 vccd1 _01927_ sky130_fd_sc_hd__nand2_1
XANTENNA__07671__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05201_ _00912_ _00913_ _00911_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__or3b_1
XFILLER_0_29_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06181_ _00649_ net132 net122 _00635_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05132_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00845_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold404 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1
+ vccd1 net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold426 _00196_ vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] vssd1 vssd1
+ vccd1 vccd1 net1106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\] vssd1 vssd1 vccd1
+ vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09940_ net461 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
X_05063_ _00792_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[2\]
+ sky130_fd_sc_hd__inv_2
Xhold459 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\] vssd1 vssd1 vccd1
+ vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09871_ net408 _01789_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__nor2_1
XANTENNA__07187__A1 _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _04168_ _04169_ net193 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08753_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
X_05965_ net212 _01656_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout182_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ _01683_ _02046_ _03259_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or3_1
X_04916_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _00656_ sky130_fd_sc_hd__inv_2
X_05896_ _01585_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__nand2_4
X_08684_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _04081_ vssd1
+ vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06698__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ net134 _01683_ _01687_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07566_ _03106_ _03116_ _03119_ _03124_ _03104_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__a221o_1
X_09305_ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06517_ net277 _02106_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__and2_2
XANTENNA__07647__C1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07497_ _01640_ _03053_ _03056_ _02390_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09236_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ _04440_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840__515 vssd1 vssd1 vccd1 vccd1 _10840__515/HI net515 sky130_fd_sc_hd__conb_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06448_ _01693_ _02047_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09167_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06379_ _01687_ _01690_ _01696_ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08118_ net759 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[8\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__mux2_1
X_09098_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04333_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ net450 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ net390 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout95_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07178__A1 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ clknet_leaf_22_wb_clk_i _00008_ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07717__A3 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07525__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10913_ net657 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06153__A2 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10844_ net519 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_67_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05699__B _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10775_ clknet_leaf_65_wb_clk_i _00596_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06147__Y _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05986__Y _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05416__A1 _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06613__B1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05416__B2 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07169__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10209_ clknet_leaf_72_wb_clk_i _00213_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08030__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05750_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__or4_1
X_05681_ net438 _01392_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07420_ net1062 _03004_ _03006_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[13\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07351_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06302_ _01967_ _01968_ net212 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05402__B _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07282_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ _00679_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09021_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04280_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__and2_1
X_06233_ _01865_ _01870_ _01880_ net114 _01882_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_135_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05896__Y _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06164_ _01820_ _01842_ _01844_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a21oi_1
Xhold201 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06073__X _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold212 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[46\]
+ vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05115_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] net447 vssd1 vssd1
+ vccd1 vccd1 _00828_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\] vssd1
+ vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__dlygate4sd3_1
X_06095_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\]
+ _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__or3_1
Xhold245 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] vssd1
+ vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08947__A_N net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold256 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _01784_ _04870_ _04901_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__o21ai_1
X_05046_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] vssd1 vssd1 vccd1 vccd1
+ _00778_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold289 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout397_A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09854_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\] _04855_ vssd1
+ vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__nand2_1
X_08805_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\] _04156_ vssd1
+ vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__nor2_1
X_09785_ _00657_ _04809_ _04808_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06383__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout185_X net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06997_ _02658_ _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08736_ net1111 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__mux2_1
XANTENNA__07064__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05948_ net253 net194 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08667_ _04076_ _04094_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__a21o_1
X_05879_ _01562_ net147 _01564_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07618_ _02208_ _03127_ _03128_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__o31a_1
X_08598_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03623_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05894__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _02838_ _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05312__B _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ clknet_leaf_0_wb_clk_i _00428_ _00065_ vssd1 vssd1 vccd1 vccd1 team_07_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07635__A2 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06127__C _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _04430_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10491_ clknet_leaf_14_wb_clk_i _00359_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07774__A1_N net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08115__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout98_X net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07571__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07874__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05885__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10827_ net502 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_7_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05997__X _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10758_ clknet_leaf_60_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[5\]
+ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06605__Y _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ clknet_leaf_34_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[21\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06053__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06920_ net174 _02511_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__and2_1
X_06851_ _02521_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05802_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\]
+ _01486_ _01487_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__and4_2
X_09570_ net482 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ _04657_ _04659_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_69_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06782_ net422 net157 _02445_ _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08521_ net858 _03982_ vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05733_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\] _00772_ _00784_
+ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08452_ _03924_ _03892_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_65_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05664_ _01256_ _01259_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_137_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] _02994_
+ net475 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__o21ai_1
X_08383_ net489 _03855_ _03858_ _03751_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__o31a_1
X_05595_ net416 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] vssd1 vssd1 vccd1
+ vccd1 _01308_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_102_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05132__B _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05628__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07265_ _02905_ _02906_ _01315_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[15\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09004_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06216_ _01850_ _01893_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__nand2_1
X_07196_ net159 _01688_ _02836_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06244__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06147_ net171 _01724_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nor2_4
XFILLER_0_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07059__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06078_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 _01765_ sky130_fd_sc_hd__nor3_1
XFILLER_0_111_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09906_ net855 net152 net150 _04891_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__a22o_1
X_05029_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05147__X _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ _04838_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] vssd1 vssd1
+ vccd1 vccd1 _04846_ sky130_fd_sc_hd__a31o_1
XANTENNA__07553__A1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _04767_ _04790_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ net931 _04132_ _04133_ vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__a21oi_1
X_09699_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] _04729_ _04742_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] vssd1 vssd1 vccd1
+ vccd1 _04747_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07522__B _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10846__521 vssd1 vssd1 vccd1 vccd1 _10846__521/HI net521 sky130_fd_sc_hd__conb_1
XANTENNA__06513__C1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05323__A _01008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10612_ clknet_leaf_40_wb_clk_i _00476_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07608__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10543_ clknet_leaf_11_wb_clk_i _00411_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05977__B net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07084__A3 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06425__Y _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10474_ clknet_leaf_27_wb_clk_i _00342_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06044__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input30_X net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10933__582 vssd1 vssd1 vccd1 vccd1 _10933__582/HI net582 sky130_fd_sc_hd__conb_1
XANTENNA__07544__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05217__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06048__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05380_ _01002_ _01023_ _01092_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_60_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05887__B _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06283__A1 _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07050_ _02692_ _02701_ _02704_ _02699_ _02703_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06001_ net132 net122 _01676_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06035__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06860__A1_N net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07952_ net269 _03346_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__or3b_1
XANTENNA__06511__B _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ _02538_ _02573_ _02536_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__o21bai_1
X_07883_ _02331_ _03291_ _03290_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__o21a_1
XANTENNA__07535__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09622_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] _04688_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_108_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06834_ _02504_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09553_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ net266 net288 net218 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a211o_1
X_06765_ _02430_ _02435_ _02436_ _02426_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_104_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08504_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ _00697_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 _03970_ sky130_fd_sc_hd__and4b_1
X_05716_ net410 _01411_ _01423_ _00826_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09484_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] vssd1
+ vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__nand2b_1
X_06696_ _02271_ _02364_ _02365_ _02367_ _02368_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_19_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05143__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08435_ net485 _03846_ _03873_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05647_ _00678_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01359_ vssd1
+ vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_121_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout148_X net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08366_ _01253_ _01381_ _03733_ _03841_ net458 vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o32a_1
X_05578_ _01289_ _01290_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07317_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ _00723_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08297_ net457 _03774_ _03694_ _00729_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07471__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ _02893_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ _02895_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06405__C _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07179_ _02822_ _02826_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__or2_1
X_10190_ clknet_leaf_80_wb_clk_i _00194_ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06702__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07774__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_4
Xfanout341 net342 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout363 net385 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
Xfanout374 net385 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
Xfanout385 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_4
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_2
XANTENNA__07533__A _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07829__A2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05988__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06436__X _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_X clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput38 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06265__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10526_ clknet_leaf_30_wb_clk_i net1010 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05994__Y _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10457_ clknet_leaf_27_wb_clk_i _00337_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07214__B1 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ clknet_leaf_4_wb_clk_i net693 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_36_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06568__A2 _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06331__B team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11009_ net638 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_74_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ _01611_ net249 _02223_ _02043_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__or4b_1
XANTENNA__08973__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05501_ net418 _00691_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ _01198_ _01213_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_16_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06481_ _01828_ _02154_ net199 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_118_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08220_ team_07_WB.instance_to_wrap.team_07.labelPixel\[0\] team_07_WB.instance_to_wrap.team_07.labelPixel\[3\]
+ team_07_WB.instance_to_wrap.team_07.labelPixel\[2\] team_07_WB.instance_to_wrap.team_07.displayPixel
+ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05432_ _01144_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XANTENNA__06346__X _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ _00717_ net470 vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__nor2_2
X_05363_ net433 _01049_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__nor2_2
XFILLER_0_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06506__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07102_ net260 _02197_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08082_ net479 _00815_ _03593_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__and3_2
XFILLER_0_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05294_ _01002_ _01006_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07033_ _01636_ net83 _02350_ _02335_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout108_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06522__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06559__A2 _02230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04253_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__or3_1
X_07935_ _03479_ _03488_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__and3b_1
XANTENNA__07508__A1 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08705__B1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_A net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07866_ _03339_ _03419_ _03420_ _03397_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09605_ _03976_ _04679_ _04680_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06817_ net270 _02487_ _02482_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_123_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07797_ _01115_ net110 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__and2_1
X_09536_ net932 net205 _04648_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__o21a_1
X_06748_ net173 _02418_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__or2_1
X_09467_ net915 net202 _04606_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__o21a_1
X_06679_ _00759_ net84 _02250_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08418_ _03655_ _03891_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07800__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09398_ net410 _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08349_ net469 _03660_ net466 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08912__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10311_ clknet_leaf_41_wb_clk_i net728 net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_105_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07087__X _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ clknet_leaf_78_wb_clk_i _00234_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06432__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ clknet_leaf_27_wb_clk_i _00183_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input38_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 net161 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
Xfanout171 _01543_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_6
Xfanout182 _01532_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10104__D team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout193 _04144_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08172__B2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06486__A1 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05230__B team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10509_ clknet_leaf_12_wb_clk_i _00377_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08033__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06342__A _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08935__A0 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06061__B _00828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05981_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\] _01633_ vssd1
+ vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__nand2_1
XANTENNA__08950__A3 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06961__A2 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _01105_ _01597_ _01604_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__and3_1
X_04932_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07651_ _03098_ _03099_ _03207_ _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__a22o_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07604__C _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06174__B1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ net174 _02013_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__nand2_1
X_07582_ _02842_ _03140_ _03118_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__o21ai_1
X_09321_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04499_ _04501_ _04503_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__o22a_1
XANTENNA__05899__Y _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06533_ _02102_ _02155_ _02153_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06464_ net274 net272 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__nor2_4
XANTENNA__06517__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\] _00730_ vssd1
+ vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05415_ _01023_ _01100_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__nor2_1
X_09183_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04396_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_32_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06395_ _01677_ _01689_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05140__B _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05346_ net190 _01000_ _01019_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__or3_2
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07977__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__B2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ net451 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05277_ _00982_ _00988_ _00989_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_116_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07016_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ _02671_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__and3_1
XANTENNA__09266__C net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08967_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] net852
+ net444 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
X_07918_ _01083_ net148 _03443_ _03441_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a31o_1
X_08898_ _04214_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\]
+ _04209_ vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07849_ net262 _03354_ _03363_ net263 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__o22a_1
XANTENNA__07901__A1 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ net535 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_79_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ net220 _04605_ net884 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a22o_1
XANTENNA__07811__A _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10791_ clknet_leaf_76_wb_clk_i _00612_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06468__A1 _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06468__B2 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08118__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06427__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__A3 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07417__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05985__B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05979__B1 _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06433__Y _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10225_ clknet_leaf_79_wb_clk_i _00229_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_7_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ clknet_leaf_15_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07705__B net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ clknet_leaf_67_wb_clk_i _00145_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload3_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10989_ net629 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_48_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06337__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05200_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00901_ vssd1 vssd1
+ vccd1 vccd1 _00913_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06180_ net286 net133 _01859_ _01860_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05131_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ _00843_ _00840_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux4_2
XFILLER_0_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold405 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\] vssd1 vssd1
+ vccd1 vccd1 net1074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold416 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\] vssd1 vssd1
+ vccd1 vccd1 net1096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold438 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] vssd1 vssd1
+ vccd1 vccd1 net1107 sky130_fd_sc_hd__dlygate4sd3_1
X_05062_ _00785_ _00789_ _00790_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__nand3_1
Xhold449 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] vssd1 vssd1
+ vccd1 vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06072__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08908__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10109__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09870_ _00827_ _01789_ net408 vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\]
+ _01448_ _04160_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_5_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06934__A2 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08752_ net1058 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
XANTENNA__07615__B _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05964_ net212 net195 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__nand2_4
X_07703_ _01686_ _01737_ _02040_ _01646_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__a2bb2o_1
X_04915_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _00655_ sky130_fd_sc_hd__inv_2
X_08683_ _04106_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04105_ vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__mux2_1
X_05895_ _01586_ _01588_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout175_A _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ net102 _02056_ _02085_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06698__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ _01704_ _02219_ _03123_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout342_A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ _04486_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06516_ _01922_ _02178_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__nor2_1
XANTENNA__07647__B1 _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ _02770_ _03054_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09235_ net227 _04441_ _04442_ net406 net958 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__a32o_1
X_06447_ _02086_ _02120_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout130_X net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04369_ _04384_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06378_ _02043_ _02050_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08117_ net799 net798 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05329_ _01008_ _01015_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__or2_1
X_09097_ net208 _04339_ _04340_ net397 net995 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06622__A1 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08048_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ net295 _03577_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout88_A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ clknet_leaf_53_wb_clk_i _00007_ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_09999_ clknet_leaf_32_wb_clk_i net1068 net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07525__B _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10912_ net656 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_98_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07541__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10843_ net518 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ clknet_leaf_66_wb_clk_i _00595_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06157__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05996__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06604__B _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06074__C1 _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06613__A1 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10208_ clknet_leaf_71_wb_clk_i _00212_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10139_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.recGen.circleDetect
+ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.circlePixel sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06129__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05680_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\] _01376_ vssd1 vssd1
+ vccd1 vccd1 _01393_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06338__Y _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10863__538 vssd1 vssd1 vccd1 vccd1 _10863__538/HI net538 sky130_fd_sc_hd__conb_1
XFILLER_0_70_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07350_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06301_ net434 _01966_ _01968_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06521__A1_N _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07281_ _02915_ _02916_ _00679_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[9\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09020_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04280_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06232_ _01670_ _01706_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06163_ net114 _01840_ _01843_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__o21a_1
Xhold202 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 _00506_ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold224 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] vssd1 vssd1
+ vccd1 vccd1 net893 sky130_fd_sc_hd__dlygate4sd3_1
X_05114_ _00826_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
Xhold235 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[43\]
+ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__dlygate4sd3_1
X_06094_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] _01776_ vssd1
+ vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold257 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\] vssd1 vssd1
+ vccd1 vccd1 net926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _01783_ net151 net727 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__o21ai_1
X_05045_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__or4bb_1
Xhold279 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\] vssd1 vssd1
+ vccd1 vccd1 net948 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09853_ _04825_ _04855_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout292_A _03033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net192 _04157_ vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__nor2_1
X_09784_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] net264 vssd1
+ vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or2_1
X_06996_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] _02649_
+ _02651_ _02659_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09306__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__mux2_1
XANTENNA__07064__C _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05947_ _01637_ _01640_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__B1 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _04080_ _04093_ _04084_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__o21ai_1
X_05878_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _01561_
+ net147 _01571_ _01559_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a32oi_2
X_07617_ _01655_ net166 _03132_ _03172_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_113_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08597_ _03623_ _04032_ net140 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07548_ _01726_ _03083_ _03085_ net201 vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o22a_1
XANTENNA__05894__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07096__B2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07479_ _01618_ _02079_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ clknet_leaf_14_wb_clk_i _00358_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09149_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07571__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ net501 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__05885__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07087__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10757_ clknet_leaf_60_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[4\]
+ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10688_ clknet_leaf_34_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[20\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06334__B _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06350__A _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ net428 _02520_ _02518_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__a21o_1
XANTENNA__08976__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05801_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] _01486_
+ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06781_ _02448_ _02452_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08520_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] vssd1 vssd1 vccd1 vccd1
+ _03983_ sky130_fd_sc_hd__and3_1
X_05732_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00772_ _00766_
+ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__a21o_1
XANTENNA__07314__A2 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08451_ net466 net473 _03640_ _03657_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_65_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05663_ _01374_ _01375_ _01346_ _01366_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__o211a_1
X_07402_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[6\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06509__B _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05413__B _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ net474 _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__nor2_1
X_05594_ _01305_ _01306_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ _00675_ _02946_ _02945_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout138_A _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05700__Y _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07264_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09003_ net247 net404 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
X_06215_ net91 _01800_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07195_ _02783_ _02832_ _02845_ _02777_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout305_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06146_ _01823_ _01826_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__or2_1
X_06077_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__nor2_1
XANTENNA__07356__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ _01779_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05028_ _00753_ _00760_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09836_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__inv_2
XANTENNA__07553__A2 _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\]
+ _02643_ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__and3_1
X_09767_ net245 _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08718_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ _04132_ net258 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__o21ai_1
X_09698_ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__inv_2
XANTENNA__07091__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08649_ _00693_ _04067_ _04059_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_25_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10885__560 vssd1 vssd1 vccd1 vccd1 _10885__560/HI net560 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_25_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10611_ clknet_leaf_40_wb_clk_i _00475_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08266__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10542_ clknet_leaf_29_wb_clk_i _00410_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06435__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ clknet_leaf_27_wb_clk_i _00341_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07777__C1 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06044__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05993__B net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11025_ net388 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07544__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__B1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10809_ clknet_leaf_67_wb_clk_i _00630_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08036__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06283__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06000_ net133 net137 net168 _01687_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07951_ net393 net110 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06902_ net430 _02106_ _00749_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07882_ _03329_ _03338_ _03409_ _03436_ _03328_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__o2111a_1
XANTENNA__07535__A2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10912__656 vssd1 vssd1 vccd1 vccd1 net656 _10912__656/LO sky130_fd_sc_hd__conb_1
X_09621_ _04666_ _04690_ _04691_ _04664_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__a32o_1
XANTENNA__07904__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] net174 vssd1 vssd1
+ vccd1 vccd1 _02504_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_108_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07940__C1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ net930 net203 _04655_ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__o21a_1
X_10869__544 vssd1 vssd1 vccd1 vccd1 _10869__544/HI net544 sky130_fd_sc_hd__conb_1
X_06764_ net99 _02417_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__xnor2_1
X_08503_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\] _03968_ vssd1 vssd1
+ vccd1 vccd1 _03969_ sky130_fd_sc_hd__nor4_1
X_05715_ net1100 _00797_ _01412_ _01426_ _01427_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a221o_1
X_09483_ net923 net203 _04615_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06695_ _02284_ _02286_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__nor2_1
XANTENNA__07342__C _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08434_ net462 _03561_ _03907_ net483 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05646_ _01357_ _01358_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_121_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08365_ net459 _03839_ _03840_ _01379_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05577_ _01282_ _01288_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07316_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ net458 _03773_ _03675_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07471__A1 _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07178_ _01665_ _01724_ _02829_ net201 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06129_ _01720_ _01735_ net283 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05785__A1 _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout320 net326 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
Xfanout342 net344 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
Xfanout353 net360 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
Xfanout364 net370 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_4
Xfanout375 net380 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_4
Xfanout386 net388 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_2
Xfanout397 net398 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_2
X_09819_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__and4_1
XANTENNA__06734__B1 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__C1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05988__B net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_10525_ clknet_leaf_28_wb_clk_i _00393_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput39 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10456_ clknet_leaf_61_wb_clk_i _00016_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07214__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10387_ clknet_leaf_4_wb_clk_i net684 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05068__X _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11008_ net387 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10981__621 vssd1 vssd1 vccd1 vccd1 _10981__621/HI net621 sky130_fd_sc_hd__conb_1
X_05500_ net418 _00691_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06480_ net143 net105 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__nor2_4
XFILLER_0_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05431_ _01077_ _01127_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05898__B _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08150_ _03635_ _03636_ vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05362_ net188 _01074_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07101_ _02754_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06506__C net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08081_ _00814_ _01429_ net229 net954 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05293_ net189 _01004_ _01005_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__nor3_1
XFILLER_0_31_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07032_ _02251_ _02686_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06661__C1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06362__X _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07177__Y _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06522__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06559__A3 _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__or2_1
XANTENNA__05138__B _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ _01084_ _03309_ _03316_ net187 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07508__A2 _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ _03359_ _03390_ _03288_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09604_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ _04678_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__nand3_1
X_06816_ _02484_ _02486_ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_123_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07796_ net276 _01115_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_123_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05154__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06747_ _02418_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__inv_2
X_09535_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ net267 _04647_ net289 net220 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__Y _03198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09466_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ net265 net288 net218 vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a211o_1
X_06678_ _02184_ _02350_ _02349_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_66_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04993__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07692__A1 _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08417_ _00717_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05629_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] _01315_
+ _01339_ _01341_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__o211ai_2
X_09397_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\] vssd1 vssd1
+ vccd1 vccd1 _04555_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08348_ _00126_ _03824_ _03801_ vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06247__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ net465 _03756_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10310_ clknet_leaf_41_wb_clk_i net747 net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09197__A1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ clknet_leaf_74_wb_clk_i net695 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06432__B net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05329__A _01008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ clknet_leaf_23_wb_clk_i _00182_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout150 _04869_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout161 _01557_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_4
Xfanout172 _01544_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
Xfanout183 _01532_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_4
XANTENNA__06707__B1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07263__B team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10965__605 vssd1 vssd1 vccd1 vccd1 _10965__605/HI net605 sky130_fd_sc_hd__conb_1
XFILLER_0_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05999__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07683__A1 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05070__Y team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05446__B1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10508_ clknet_leaf_12_wb_clk_i _00376_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ clknet_leaf_42_wb_clk_i _00323_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07199__B1 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06342__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06577__B1_N _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05980_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] _01633_ _01641_
+ _01660_ _01673_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\]
+ sky130_fd_sc_hd__a2111oi_2
XTAP_TAPCELL_ROW_72_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04931_ net422 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10088__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ net250 _01734_ _02371_ _03114_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06174__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06174__B2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06601_ net123 _01652_ _02014_ net156 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a211o_1
XANTENNA__07910__A2 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ net130 net138 _01719_ _01903_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a31o_1
X_09320_ _00661_ _04500_ net225 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06532_ _02188_ _02199_ _02205_ _02183_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or4b_1
XANTENNA__06357__X _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04449_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06463_ _02053_ _02136_ _02135_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06517__B _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08202_ net460 _01383_ _03680_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05414_ net433 _01062_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ net207 _04401_ _04402_ net403 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_32_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06394_ _01693_ _01696_ _02052_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08133_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ _03619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05345_ net433 _01048_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout120_A _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08064_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net391 net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ _03585_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05276_ net422 _00983_ _00670_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07015_ _02671_ vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10918__662 vssd1 vssd1 vccd1 vccd1 net662 _10918__662/LO sky130_fd_sc_hd__conb_1
X_08966_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] net748
+ net444 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07917_ net272 _03354_ _03363_ net269 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__o22a_1
X_08897_ _00708_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ net479 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07848_ _01679_ _03380_ _03388_ _01689_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o22a_1
XANTENNA__07901__A2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ net431 net110 _03275_ _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_116_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ net884 net204 _04636_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__o21a_1
XANTENNA__07811__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10790_ clknet_leaf_76_wb_clk_i _00611_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07665__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09449_ _01415_ _04589_ _04586_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a21o_1
XANTENNA__08862__B1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06427__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07968__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05979__A1 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10224_ clknet_leaf_72_wb_clk_i _00228_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ clknet_leaf_15_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ clknet_leaf_67_wb_clk_i _00144_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07561__X _03120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10988_ net628 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_128_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06337__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05130_ _00835_ _00841_ _00842_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07959__A2 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08044__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] vssd1 vssd1 vccd1
+ vccd1 net1075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold428 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] vssd1 vssd1
+ vccd1 vccd1 net1097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold439 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__dlygate4sd3_1
X_05061_ _00790_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] _01448_
+ _04160_ net862 vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_110_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08751_ net1146 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__mux2_1
X_05963_ net215 net196 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07702_ net86 _01635_ _03257_ _03255_ _03251_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__o311a_1
X_04914_ net971 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
X_05894_ _01574_ _01575_ _00715_ _01569_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a211oi_2
X_08682_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04082_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07633_ _01660_ _02167_ _03080_ _03117_ _03190_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a41o_1
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07564_ net102 _03078_ _03121_ _03122_ _01646_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ _04486_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a21o_1
X_06515_ _02054_ _02115_ _02155_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07647__A1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ _00685_ _00941_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09234_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04435_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__a21o_1
X_06446_ net167 _02069_ _02088_ _02110_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a211o_1
XANTENNA__05151__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04384_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06377_ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout123_X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08116_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\] net806
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1 vssd1 vccd1 vccd1
+ _00116_ sky130_fd_sc_hd__mux2_1
X_05328_ _01008_ _01015_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__nor2_1
X_09096_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ _04337_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08047_ net450 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ net390 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05259_ _00671_ net424 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10253__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__04989__Y _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06386__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07806__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ clknet_leaf_33_wb_clk_i _00001_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07583__B1 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ net491 _04241_ vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07822__A _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ net655 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07541__B _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ net517 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__06438__A _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10773_ clknet_leaf_65_wb_clk_i _00594_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05996__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10207_ clknet_leaf_72_wb_clk_i _00211_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.borderGen.synchronized_rectangle_pixel
+ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06129__A1 _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ clknet_leaf_48_wb_clk_i _00127_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09866__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07451__B net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08039__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06300_ net184 _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07280_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06231_ _01892_ _01895_ _01896_ _01909_ _01889_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a41o_1
XFILLER_0_116_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10904__569 vssd1 vssd1 vccd1 vccd1 _10904__569/HI net569 sky130_fd_sc_hd__conb_1
XANTENNA__06852__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10276__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06162_ net120 _01797_ _01804_ _01840_ net113 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a32o_1
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] vssd1 vssd1
+ vccd1 vccd1 net872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold214 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__dlygate4sd3_1
X_05113_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\] vssd1 vssd1 vccd1
+ vccd1 _00826_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_113_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold225 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__dlygate4sd3_1
X_06093_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\]
+ _01775_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold236 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _00467_ vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _01783_ _04870_ _04900_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__o21ai_1
X_05044_ _00652_ _00775_ _00763_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07907__A _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09852_ net264 _04854_ _04856_ net243 net1064 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__a32o_1
X_08803_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\] _04156_ vssd1
+ vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__xor2_1
X_09783_ net264 _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand2b_2
X_06995_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] _02650_
+ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__nor2_1
X_08734_ net1125 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05946_ net98 net88 net271 _01638_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a31o_1
X_05877_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01555_
+ _01546_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08665_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04047_ _04072_ _04089_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o311a_1
X_07616_ net125 _01676_ _03173_ _02262_ net165 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a32o_1
XANTENNA__06258__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\] _03621_
+ net848 vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__o31ai_1
XANTENNA__05162__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ _03105_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07096__A2 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ _01626_ _01635_ _02176_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__or3b_1
XANTENNA__08293__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ net227 _04428_ _04429_ net406 net1009 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_20_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06429_ _01722_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07089__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ net206 _04377_ _04378_ net401 net1020 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__a32o_1
XANTENNA__09242__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10769__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06056__B1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09079_ net208 _04326_ _04327_ net400 net985 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06280__X _01957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07817__A _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10008__SET_B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__B1 _02930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ net500 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10756_ clknet_leaf_61_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\]
+ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06455__X _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10687_ clknet_leaf_34_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[19\]
+ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_93_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06631__A _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06350__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830__505 vssd1 vssd1 vccd1 vccd1 _10830__505/HI net505 sky130_fd_sc_hd__conb_1
X_05800_ _01490_ _01493_ _01491_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__and4bb_1
X_06780_ _00984_ net173 _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05731_ _00709_ _00710_ _01436_ _01434_ net486 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a32o_1
XFILLER_0_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05253__Y _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08450_ _03662_ _03815_ _03922_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__o211a_1
X_05662_ _01255_ _01257_ _01278_ _01323_ _00679_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_106_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07401_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\] _02992_
+ net476 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06509__C _02042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08381_ _03856_ team_07_WB.instance_to_wrap.team_07.defusedGen.defusedPixel team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05593_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] vssd1 vssd1 vccd1
+ vccd1 _01306_ sky130_fd_sc_hd__or3b_2
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07332_ net426 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07263_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06214_ _01807_ _01892_ _01893_ _01820_ _01891_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a221o_1
X_09002_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ net2 _04252_ _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_60_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07194_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06145_ net91 _01803_ _01825_ net101 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout200_A _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06076_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] vssd1 vssd1 vccd1
+ vccd1 _01763_ sky130_fd_sc_hd__and3b_1
XFILLER_0_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] _01778_
+ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05027_ net282 _00751_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__nor2_1
XANTENNA_input5_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ _04840_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__and3_1
X_09766_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] _04790_ _04767_
+ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a21boi_1
X_06978_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _02643_
+ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__xor2_1
X_08717_ _04128_ _04130_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__nor2_1
X_05929_ net281 net270 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09697_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ net246 _04742_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__and4_1
XANTENNA__06259__Y _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ _04054_ _04075_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a21o_1
XANTENNA__06513__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08579_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ _03618_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10610_ clknet_leaf_40_wb_clk_i net887 net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10541_ clknet_leaf_30_wb_clk_i _00409_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10472_ clknet_leaf_27_wb_clk_i _00340_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06029__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07777__B1 _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07529__B1 _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11024_ net643 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08378__A _00711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10808_ clknet_leaf_76_wb_clk_i _00629_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10739_ clknet_leaf_62_wb_clk_i _00569_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09937__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07950_ _03471_ _03472_ _03503_ _03504_ _03502_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06901_ _02527_ _02542_ _02570_ _02571_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
X_07881_ _03417_ _03418_ _03434_ _03435_ _03412_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09620_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] _04688_ vssd1
+ vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__nand2_1
XANTENNA__07535__A3 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ _02501_ _02502_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09551_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ net266 net287 net218 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a211o_1
X_06763_ _02425_ _02431_ _02434_ _02423_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08502_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__or4b_1
X_05714_ net410 _00827_ _01423_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__nor3_1
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09482_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ net266 _04612_ _04614_ net218 vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a221o_1
X_06694_ _01624_ net84 _02313_ net249 _02366_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08433_ net462 _03857_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05645_ net415 _00676_ _00677_ _01356_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__o31a_1
XFILLER_0_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08248__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05711__Y _01424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08364_ _03678_ _03731_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__or2_1
X_05576_ _01282_ _01288_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05440__A _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08295_ net415 _03678_ _03772_ net459 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07246_ _00720_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ _02894_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07177_ net201 _02828_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__nand2_2
X_06128_ net286 net107 _01691_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__or3_1
XFILLER_0_112_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06271__A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06059_ net1123 _01633_ _01746_ _01747_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\]
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_111_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout310 net315 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05785__A2 _01481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_4
Xfanout332 net351 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_4
Xfanout343 net344 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
Xfanout354 net360 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_4
Xfanout365 net370 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 net380 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
X_09818_ net1149 _04830_ _04831_ _04832_ vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__o22a_1
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_2
Xfanout398 net399 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07814__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09749_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] _04777_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07533__C _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08487__A1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput18 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10524_ clknet_leaf_13_wb_clk_i _00392_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ sky130_fd_sc_hd__dfrtp_1
Xinput29 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10015__RESET_B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06670__B1 _02027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10455_ clknet_leaf_61_wb_clk_i _00015_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10386_ clknet_leaf_4_wb_clk_i net683 net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05509__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11007_ net387 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06725__B2 _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05244__B _00956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05430_ _01026_ _01110_ _01106_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05898__C _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06356__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05361_ _01005_ _01019_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06075__B _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ _02726_ _02729_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__and2b_1
X_08080_ _03591_ _03592_ _00815_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07453__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05292_ _00675_ _00998_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07031_ net260 net83 _02335_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a21o_1
XANTENNA__05464__A1 _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05464__B2 _01112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09386__B _01424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08402__A1 _00711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10836__511 vssd1 vssd1 vccd1 vccd1 _10836__511/HI net511 sky130_fd_sc_hd__conb_1
XANTENNA__06413__B1 _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08982_ _00664_ _04249_ _04250_ _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ _03305_ _03442_ _03444_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07864_ _03352_ _03360_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06716__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] _04678_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06815_ net282 net430 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_123_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ _03348_ _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__nand2b_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05154__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _00666_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] vssd1 vssd1
+ vccd1 vccd1 _04647_ sky130_fd_sc_hd__a21oi_1
X_06746_ _00670_ _00983_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ net218 _04605_ net937 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07141__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06677_ _01636_ net84 _02250_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08416_ net465 net468 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05628_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] net439
+ net441 _01338_ _01340_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__o311a_1
X_09396_ net410 net413 _01475_ _04554_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08347_ _03753_ _03814_ _03818_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05559_ _01269_ _01271_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _03638_ _03641_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07229_ _02860_ _02856_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10240_ clknet_leaf_74_wb_clk_i net687 net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06404__B1 _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ clknet_leaf_27_wb_clk_i _00181_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout140 _03625_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout151 net153 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_2
Xfanout173 _01544_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_4
Xfanout195 _01518_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05064__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05999__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05351__Y _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07683__A2 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10507_ clknet_leaf_12_wb_clk_i _00375_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07719__B _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07772__A1_N _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10438_ clknet_leaf_42_wb_clk_i _00322_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07199__A1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ clknet_leaf_3_wb_clk_i net671 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07735__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04930_ net421 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XANTENNA__09950__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06174__A2 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ _01804_ _02013_ net251 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a21o_1
X_07580_ _03136_ _03138_ _03129_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05921__A2 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06531_ _01624_ _02166_ net84 _02204_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_0_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04449_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__a21o_1
X_06462_ net104 net164 _02104_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07674__A2 _02282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08201_ net416 net460 _01257_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__and3b_1
X_05413_ _01047_ _01109_ _01121_ _01125_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__and4b_1
X_09181_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06393_ _00649_ _02065_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_32_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05344_ _00668_ _01056_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__nor2_4
X_08132_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ _03618_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08063_ net453 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__and2b_1
X_05275_ _00979_ _00987_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__nand2_2
XFILLER_0_109_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout113_A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07014_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck
+ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__and2b_2
XFILLER_0_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08387__B1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07916__Y _03471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08965_ net417 net750 net444 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout482_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _03455_ _03461_ _03466_ _03470_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__a22oi_2
X_10988__628 vssd1 vssd1 vccd1 vccd1 _10988__628/HI net628 sky130_fd_sc_hd__conb_1
X_08896_ _04213_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ _04209_ vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__mux2_1
XANTENNA__05165__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ net269 _03392_ _03401_ _03398_ _03393_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07778_ net431 net110 _03330_ _03332_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__o211a_1
X_09517_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ net267 net289 net221 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06729_ _02079_ _02149_ net83 _02066_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09448_ net925 net202 _04594_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__o21a_1
XANTENNA__07665__A2 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09379_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04541_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05979__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10223_ clknet_leaf_79_wb_clk_i _00227_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06928__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ clknet_leaf_15_wb_clk_i net846 net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10085_ clknet_leaf_67_wb_clk_i _00143_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold7 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10987_ net627 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_58_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05081__Y team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07449__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__A3 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold407 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] vssd1 vssd1
+ vccd1 vccd1 net1076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold418 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 net1087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09945__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05060_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] _00788_ vssd1
+ vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__nand2_1
Xhold429 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] vssd1 vssd1
+ vccd1 vccd1 net1098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07041__B1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08750_ net1039 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__mux2_1
X_05962_ net196 _01645_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07701_ net112 _01921_ _02176_ _02332_ _02216_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__a221o_1
X_04913_ net860 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_08681_ _04034_ _04083_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05893_ _01586_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__inv_2
X_07632_ _01632_ _02182_ _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__and3b_1
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05713__A _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ _01543_ _01701_ _02743_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ net225 _04488_ _04489_ net396 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06514_ _01711_ _02047_ _02184_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a31o_1
X_07494_ net277 _00749_ net118 net89 vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__a31o_1
XANTENNA__07647__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06445_ net275 net279 net263 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__or3_4
XFILLER_0_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout328_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09164_ net1124 net403 net206 _04389_ vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__a22o_1
X_06376_ _02047_ _02049_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__and2_2
XFILLER_0_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08115_ net770 net765 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05327_ _01039_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
X_09095_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ _04337_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout116_X net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08046_ _03576_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ net454 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__mux2_1
X_05258_ net422 _00672_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05189_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00901_ vssd1 vssd1
+ vccd1 vccd1 _00902_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ clknet_leaf_32_wb_clk_i _00018_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06386__A2 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A1 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08948_ _00709_ net414 _04234_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared
+ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a31o_1
XFILLER_0_99_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08879_ _01109_ _04198_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a21oi_1
X_10910_ net654 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XANTENNA__07822__B net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ net516 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__06438__B _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10772_ clknet_leaf_66_wb_clk_i _00593_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07638__A2 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06454__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06460__Y _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10206_ clknet_leaf_71_wb_clk_i _00210_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07574__A1 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07574__B2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ clknet_leaf_53_wb_clk_i team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ clknet_leaf_46_wb_clk_i _00126_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ sky130_fd_sc_hd__dfxtp_4
XANTENNA__06129__A2 _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06629__A _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05252__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06230_ _01821_ _01890_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06161_ net113 _01840_ _01841_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07894__S net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold204 team_07_WB.instance_to_wrap.ssdec_sck vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__dlygate4sd3_1
X_05112_ net951 _00817_ _00823_ net1005 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold215 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[30\]
+ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__dlygate4sd3_1
X_06092_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] _01774_ vssd1
+ vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__or2_1
Xhold226 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[40\]
+ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold248 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _01782_ net151 net737 vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o21ai_1
X_05043_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\]
+ _00773_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__and3_1
Xhold259 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07907__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__inv_2
X_08802_ _04155_ _04156_ net193 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__a21oi_1
X_09782_ _00655_ _00656_ _00764_ _04806_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a41o_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06994_ _02652_ _02657_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__nand2_1
XANTENNA__06773__C1 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ net1152 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ net233 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__mux2_1
X_05945_ net98 net89 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout180_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ _04085_ _04090_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a22oi_2
X_05876_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] _01561_
+ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__nand2_2
XANTENNA__07868__A2 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07615_ _02873_ _03120_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__nand2_1
XANTENNA__08457__C _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08595_ _03622_ _04031_ net145 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__o21a_1
XANTENNA__06258__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05162__B _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ _02235_ _02734_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07477_ net261 _01619_ _02779_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09216_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06428_ _01722_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06359_ _01689_ _01936_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__nor2_2
XANTENNA__07089__B _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06056__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09078_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ net409 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ net291 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a221o_1
XANTENNA__07817__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout93_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07556__A1 _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05353__A _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ net499 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XANTENNA__05072__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06736__X team_07_WB.instance_to_wrap.team_07.recHEART.heartDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ clknet_leaf_61_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[2\]
+ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10686_ clknet_leaf_34_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[18\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10207__Q team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08744__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06350__C net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__RESET_B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05730_ _00711_ _01435_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06359__A _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05263__A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05661_ _01300_ _01373_ _01278_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07400_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ _02990_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06509__D _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08380_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.boomGen.boomPixel vssd1 vssd1 vccd1 vccd1 _03856_
+ sky130_fd_sc_hd__and2_1
X_05592_ net417 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] vssd1 vssd1 vccd1
+ vccd1 _01305_ sky130_fd_sc_hd__or3b_2
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07331_ _00965_ _01175_ _01190_ _01192_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07262_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08861__X _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ net2 net362 vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06213_ _01805_ _01807_ _01890_ _01892_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_104_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09676__Y _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07193_ _02822_ _02826_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06144_ _01802_ _01824_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06822__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06075_ _01748_ _01761_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ net837 net152 net150 _04889_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__a22o_1
X_05026_ net260 _00759_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout395_A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05157__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ net264 _04842_ _04843_ net243 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09765_ _04767_ _04791_ _04792_ net245 net1019 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a32o_1
X_06977_ _02643_ _02644_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout183_X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06761__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ _04131_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ _04128_ vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__mux2_1
X_05928_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net285
+ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__or2_1
X_09696_ _00700_ _04730_ _04743_ _04744_ _04734_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__o311a_1
XFILLER_0_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08647_ _04058_ _04060_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__and3b_1
X_05859_ _01548_ _01550_ _01551_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _03997_ _04022_ _03996_ vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07529_ net168 net104 _02110_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ clknet_leaf_30_wb_clk_i _00408_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10471_ clknet_leaf_27_wb_clk_i _00339_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10365__SET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06029__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout96_X net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05348__A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10853__528 vssd1 vssd1 vccd1 vccd1 _10853__528/HI net528 sky130_fd_sc_hd__conb_1
XANTENNA__07266__C team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11023_ net388 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05067__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07563__A _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05960__B1 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07162__C1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07701__B2 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05370__X _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ clknet_leaf_70_wb_clk_i _00628_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ clknet_leaf_57_wb_clk_i _00568_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10669_ clknet_leaf_26_wb_clk_i net944 net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08841__B _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08965__A0 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10644__RESET_B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06440__A1 _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ _00746_ _02568_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__or2_1
X_07880_ net106 _03381_ _03387_ _01692_ _03380_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o32a_1
XFILLER_0_37_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09390__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06831_ net160 _02500_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09550_ net888 net203 _04654_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ _02424_ _02425_ _02433_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nor3_1
X_08501_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] _00657_ vssd1 vssd1
+ vccd1 vccd1 _03967_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05713_ _01413_ _01424_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__nor2_1
X_09481_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04613_ net290 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o21a_1
X_06693_ _02209_ _02259_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08432_ _03631_ _03637_ _03901_ _03905_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_19_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05644_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] _01356_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ _01256_ _03729_ _03838_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05575_ _01286_ _01287_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06657__A1_N _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07314_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ _00722_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ sky130_fd_sc_hd__a31oi_1
X_08294_ net460 _03771_ _03680_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_116_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07245_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout310_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _00807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07208__B1 _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07176_ net185 _01901_ net196 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07759__A1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06127_ net283 _01720_ _01735_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10956__596 vssd1 vssd1 vccd1 vccd1 _10956__596/HI net596 sky130_fd_sc_hd__conb_1
X_06058_ _01641_ _01738_ _01744_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__or3_1
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 net313 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05009_ net42 net40 net43 _00744_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__and4_1
Xfanout322 net326 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
Xfanout333 net337 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout344 net350 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_4
Xfanout355 net360 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
Xfanout366 net369 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
Xfanout377 net379 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
X_09817_ _00657_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] vssd1
+ vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__nor2_1
Xfanout388 net75 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_2
Xfanout399 _00807_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09748_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ _04777_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__nand3_1
XFILLER_0_69_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _04704_ vssd1
+ vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_66_wb_clk_i_X clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10523_ clknet_leaf_12_wb_clk_i _00391_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput19 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06670__A1 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_row
+ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10385_ clknet_leaf_4_wb_clk_i net694 net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06973__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11006_ net386 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07686__B1 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05697__C1 _00962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06356__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09948__A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05360_ net190 _01004_ _01010_ _01071_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05291_ _00993_ _00995_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__or2_4
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07030_ net128 _01677_ _01708_ _02684_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06661__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05464__A2 _01103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06661__B2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10875__550 vssd1 vssd1 vccd1 vccd1 _10875__550/HI net550 sky130_fd_sc_hd__conb_1
XANTENNA__06413__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__nand3_1
XANTENNA__05419__C _01039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ _03311_ _03324_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07863_ net107 _03321_ _03326_ _01692_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07913__A1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06716__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ net1107 _04678_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__xor2_1
X_06814_ net276 net430 _02484_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07794_ net277 _01069_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07490__X _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09533_ net907 net205 _04646_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__o21a_1
X_06745_ _00673_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ _02409_ _02416_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ net217 _04605_ net874 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__a22o_1
XANTENNA__07677__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06676_ _01639_ _02348_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08415_ _03646_ _03889_ _03657_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__a21oi_1
X_05627_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] _01319_
+ _01328_ net417 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__o22a_1
X_09395_ _01425_ _04551_ _04553_ _02984_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout146_X net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08346_ _03657_ _03820_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05558_ _01254_ _01268_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08277_ net468 _00717_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__nor2_1
X_05489_ _00688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07228_ _02081_ _02775_ _02877_ _02878_ _02767_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__a32o_1
XANTENNA__06652__A1 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06282__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07159_ _02065_ net81 _02736_ _02807_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10170_ clknet_leaf_27_wb_clk_i _00180_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout130 _01577_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_4
XFILLER_0_100_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout141 net142 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
Xfanout163 _02745_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 net175 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_4
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06707__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 net198 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_4
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07668__B1 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__B _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06340__B1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07683__A3 _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07559__Y _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06643__A1 _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10506_ clknet_leaf_15_wb_clk_i _00374_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06192__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10859__534 vssd1 vssd1 vccd1 vccd1 _10859__534/HI net534 sky130_fd_sc_hd__conb_1
XANTENNA__07719__C _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10437_ clknet_leaf_42_wb_clk_i _00321_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07199__A2 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ clknet_leaf_5_wb_clk_i net717 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06920__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10299_ clknet_leaf_24_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[12\]
+ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06530_ _02202_ _02203_ _01618_ _02164_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07659__B1 _02835_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06367__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07123__A2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06461_ _00747_ _00755_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__or2_2
XFILLER_0_34_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08200_ net415 _03678_ _03677_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__o21ai_1
X_05412_ _01054_ _01117_ _01122_ _01124_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__and4b_1
X_09180_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06392_ net282 net279 _01621_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__and3_2
XANTENNA__06654__X _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05421__D _01103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08131_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__or2_1
X_05343_ net433 _00669_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__nand2_4
XFILLER_0_71_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06373__Y _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ net1053 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ net295 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__mux2_1
X_05274_ net421 _00984_ _00983_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07013_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle
+ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08387__A1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06830__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08964_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] net796
+ net444 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
X_07915_ net252 _03376_ _03469_ _03468_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__a31o_1
X_08895_ _00708_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ net479 vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05165__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _03345_ _03395_ _03399_ _03400_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07661__A _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _00669_ net120 _02212_ _01104_ _02191_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a221o_1
XANTENNA__06570__B1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04989_ net464 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09516_ net901 net204 _04635_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__o21a_1
X_06728_ net261 _02149_ net83 _02134_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_91_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ net265 _04593_ net287 net217 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06659_ net273 _02331_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09378_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04541_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ net459 _03727_ _03728_ _03732_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__o31a_1
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06724__B _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10222_ clknet_leaf_73_wb_clk_i _00226_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_10971__611 vssd1 vssd1 vccd1 vccd1 _10971__611/HI net611 sky130_fd_sc_hd__conb_1
XFILLER_0_101_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07050__A1 _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ clknet_leaf_15_wb_clk_i net715 net323 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07050__B2 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ clknet_leaf_67_wb_clk_i _00142_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09770__B _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10986_ net626 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_128_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10488__RESET_B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08853__A2 _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06915__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07813__B1 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold408 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold419 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\] vssd1 vssd1
+ vccd1 vccd1 net1088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07041__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05961_ net126 _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__nor2_4
XFILLER_0_40_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07700_ net260 _01627_ _02150_ _03250_ _03252_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__o311a_1
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_04912_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _00652_ sky130_fd_sc_hd__inv_2
X_08680_ _04103_ _04104_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__a21o_1
X_05892_ _01561_ _01568_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__xor2_2
XFILLER_0_24_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07631_ _01708_ _02263_ _03188_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07481__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06368__Y _02042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _01740_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__nor2_1
XANTENNA__05713__B _01424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ _04486_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__or2_1
X_06513_ net87 net85 _02186_ _01660_ _02079_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__o2111a_1
X_07493_ _02128_ net83 _03052_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09232_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04435_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__and3_1
X_06444_ _02084_ _02114_ _02117_ _02109_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__o31a_1
XFILLER_0_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09163_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ _04388_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_118_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06375_ net186 net178 _02048_ _01684_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08114_ net755 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[4\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__mux2_1
X_05326_ net424 _00984_ _00985_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__o21a_1
X_09094_ net208 _04336_ _04338_ net397 net1046 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08045_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ net450 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__mux2_1
X_05257_ net431 net393 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__nand2_2
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout109_X net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05188_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ _00899_ _00900_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux4_2
XFILLER_0_12_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09996_ clknet_leaf_32_wb_clk_i _00035_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09871__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ net491 _04240_ vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10232__D net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _04199_ _04200_ _04202_ _00964_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__o31a_1
XFILLER_0_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07829_ _01058_ net214 net195 _01095_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a22o_1
X_10840_ net515 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05897__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ clknet_leaf_66_wb_clk_i _00592_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10581__RESET_B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821__496 vssd1 vssd1 vccd1 vccd1 _10821__496/HI net496 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_91_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10205_ clknet_leaf_81_wb_clk_i _00209_ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07574__A2 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__A team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.recMOD.modSquaresDetect
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel
+ sky130_fd_sc_hd__dfrtp_1
X_10067_ clknet_leaf_46_wb_clk_i _00125_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.frameBufferLowNibble
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload1_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10969_ net609 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06364__B _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06160_ net113 _01840_ _01807_ _01805_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08860__A _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05111_ net1101 _00824_ _00825_ net1005 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold205 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[6\]
+ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06091_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ _01773_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_113_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold216 _00490_ vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _00500_ vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__dlygate4sd3_1
X_05042_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] _00773_ vssd1
+ vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__nand2_1
Xhold249 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08071__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ _04850_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__and3_1
X_11015__640 vssd1 vssd1 vccd1 vccd1 _11015__640/HI net640 sky130_fd_sc_hd__conb_1
XFILLER_0_42_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08801_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] _04154_ vssd1
+ vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__or2_1
X_06993_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _02651_
+ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__or2_1
X_09781_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] _00654_ vssd1
+ vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__nand2_1
XANTENNA__06773__B1 _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08732_ net982 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
X_05944_ net96 net93 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__nor2_1
XANTENNA__09711__B1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ _04049_ _04050_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ _04086_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__o221a_1
X_05875_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] net146
+ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout173_A _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__A3 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07614_ net104 net162 _03134_ _03171_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__a211o_1
XANTENNA__05879__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10339__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08594_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03621_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07545_ _03098_ _03099_ _03103_ _02055_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout340_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07476_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sck
+ sky130_fd_sc_hd__and2_1
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09215_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06427_ net275 net279 _00045_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09146_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06358_ _02031_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06056__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05309_ _01021_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09077_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06289_ net437 net131 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06561__Y _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ net451 net448 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout86_A _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ clknet_leaf_79_wb_clk_i _00084_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07325__S _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10762__RESET_B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06531__A3 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05921__X _01615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ net498 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06819__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10754_ clknet_leaf_62_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10685_ clknet_leaf_26_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[17\]
+ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06184__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10137__D team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06350__D _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10119_ clknet_leaf_45_wb_clk_i _00157_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06359__B _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05660_ _01369_ _01372_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__nor2_1
XANTENNA__05263__B net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05591_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] vssd1 vssd1 vccd1
+ vccd1 _01304_ sky130_fd_sc_hd__or3b_2
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ _02942_ _02944_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07483__A1 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07261_ _00718_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ _02903_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09000_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ net1 _04268_ vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06212_ net109 _01801_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__nand2_1
X_07192_ _02830_ _02833_ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06143_ net215 _01799_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06074_ _01395_ _01408_ _01759_ _01760_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__o211a_1
X_09902_ _01778_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__nand2_1
X_05025_ net278 _00753_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__or2_2
XFILLER_0_111_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09833_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\] _04840_ vssd1
+ vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09764_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\]
+ _04783_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 _04792_ sky130_fd_sc_hd__a31o_1
X_06976_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _02641_
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__nor2_1
XANTENNA__09571__D _01421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08715_ net259 _01756_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__and3_1
X_05927_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net285
+ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__nor2_4
X_09695_ net246 _04742_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout176_X net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05858_ _01550_ _01551_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__nand2_1
X_08646_ _01475_ _01480_ _04070_ net478 vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07710__A2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10102__RESET_B net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05789_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col
+ _01436_ _01434_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a32o_1
X_08577_ _03618_ _04021_ net140 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06556__Y _02230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ net102 _03079_ _03082_ net155 vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07459_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net391 net293 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ _03030_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[7\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10470_ clknet_leaf_11_wb_clk_i _00338_ net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06029__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ net323 _04358_ net1025 vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__a41o_1
XANTENNA__07777__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05788__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07529__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11022_ net388 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout89_X net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05916__X _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07934__C1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05960__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07162__B1 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07701__A2 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ clknet_leaf_70_wb_clk_i _00627_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07465__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10737_ clknet_leaf_57_wb_clk_i _00567_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10668_ clknet_leaf_26_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[0\]
+ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07217__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10599_ clknet_leaf_34_wb_clk_i _00463_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06728__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06830_ net159 _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07940__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ _00973_ net198 _02430_ _02432_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a211o_1
X_08500_ _00656_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__nor2_1
X_05712_ _01424_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06692_ net175 _01722_ _02014_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a21oi_2
X_09480_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\] vssd1
+ vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08431_ _03663_ _03903_ _03904_ _00703_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a221o_1
X_05643_ _01354_ _01355_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _00730_ _01258_ _03725_ _03837_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o31a_1
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05574_ _01284_ _01285_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07313_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[1\]
+ sky130_fd_sc_hd__and2b_1
X_08293_ net417 _00730_ _01258_ _03687_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__o31a_1
XFILLER_0_73_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07244_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06392__X _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07175_ _02822_ _02826_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06126_ _01797_ _01804_ net117 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07759__A2 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06057_ _01644_ _01739_ _01741_ _01745_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout301 net327 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
X_05008_ net387 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_4
Xfanout323 net325 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_4
Xfanout334 net336 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
Xfanout345 net347 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
Xfanout356 net358 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
Xfanout367 net369 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_2
X_09816_ _04829_ _04831_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__and2_1
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07392__B1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _04779_ _04778_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06959_ _02608_ _02611_ _02629_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09678_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\] net246 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08495__A _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07695__A1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ _04051_ _04056_ _00707_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_64_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10522_ clknet_leaf_12_wb_clk_i _00390_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10453_ clknet_leaf_21_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_col
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05359__A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10384_ clknet_leaf_3_wb_clk_i net675 net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11005_ net386 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05365__Y _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05290_ _00988_ _00989_ _00982_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06661__A2 _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06372__B _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06413__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__nand4_1
XFILLER_0_11_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07931_ _03314_ _03484_ _03485_ net252 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07862_ net272 _03414_ _03416_ net270 vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__o22a_1
X_09601_ _04677_ _04678_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__nor2_1
XANTENNA__06716__A3 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06813_ _02479_ _02481_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__nand2_1
X_07793_ net278 _01069_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09532_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ net267 _04638_ _04645_ net220 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a221o_1
X_06744_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ _02415_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__nand2_1
XANTENNA__06387__X _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09463_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00820_ net265 vssd1 vssd1
+ vccd1 vccd1 _04605_ sky130_fd_sc_hd__and3_4
XANTENNA__07677__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ net96 _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout253_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06547__B net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08414_ net472 _03643_ _03815_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05626_ net416 _00679_ _01327_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09394_ net413 _01416_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08345_ _03631_ _03662_ _03821_ _03659_ _03629_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o221a_1
X_05557_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] vssd1 vssd1 vccd1
+ vccd1 _01270_ sky130_fd_sc_hd__or3_2
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08276_ net129 _03670_ _03754_ _03654_ vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__a31o_1
X_05488_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07227_ net251 _01655_ _02276_ _02877_ _02040_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10256__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ _02060_ _02112_ _02810_ _02809_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a31o_1
XANTENNA__09051__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06109_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ _01791_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__nor3_1
X_07089_ net253 _01658_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05907__A _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout120 _01607_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_4
Xfanout131 _01577_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_4
Xfanout142 _01697_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_4
Xfanout153 _04868_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout164 _02055_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_4
Xfanout175 _01544_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_4
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_83_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05913__Y _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07668__A1 _02081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06340__A1 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06340__B2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07569__A _01611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ clknet_leaf_15_wb_clk_i _00373_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06192__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ clknet_leaf_42_wb_clk_i _00320_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10367_ clknet_leaf_5_wb_clk_i net676 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10298_ clknet_leaf_50_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[11\]
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07659__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06367__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06460_ net262 _00755_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__nor2_4
XFILLER_0_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05411_ net191 _01015_ _01043_ _01114_ _01123_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06391_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] _00755_
+ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_32_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08130_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05342_ net433 _00669_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__and2_2
XFILLER_0_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ net1033 net1177 net295 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__mux2_1
X_05273_ _00985_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ _02663_ _02662_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06670__X _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08963_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] net793
+ net444 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
X_07914_ _01689_ _03381_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__nor2_1
X_08894_ _04212_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ _04209_ vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
XANTENNA__07347__B1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07845_ _01077_ net110 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout370_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ _00669_ net118 vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__nand2_1
X_04988_ team_07_WB.instance_to_wrap.audio vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
X_09515_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ net268 net290 net221 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__a211o_1
X_06727_ _02395_ _02396_ _02399_ _01639_ _01630_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06277__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09446_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ net413 _04585_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__or3b_1
X_06658_ net284 net269 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05609_ net442 net441 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__nor2_1
X_10925__669 vssd1 vssd1 vccd1 vccd1 net669 _10925__669/LO sky130_fd_sc_hd__conb_1
X_09377_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04538_ _04540_ _04542_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__o22a_1
X_06589_ net123 _01654_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08328_ _00683_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ _03804_ _03747_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08259_ net487 _00727_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06580__X _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10221_ clknet_leaf_78_wb_clk_i _00225_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06740__B _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__S _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ clknet_leaf_16_wb_clk_i net698 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ clknet_leaf_67_wb_clk_i _00141_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06010__B1 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05372__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10985_ net625 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10826__501 vssd1 vssd1 vccd1 vccd1 _10826__501/HI net501 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_48_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07510__B1 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07813__A1 _01112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07813__B2 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold409 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06490__X _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ clknet_leaf_56_wb_clk_i _00310_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07041__A2 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05960_ _01574_ _01575_ _01649_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a21o_4
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04911_ net478 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05891_ _01579_ _01581_ _01584_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__and3_2
XFILLER_0_45_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07630_ _02070_ _03120_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07561_ net169 _02744_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__or2_2
X_09300_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ _04486_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nand2_1
X_06512_ _02120_ _02185_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07492_ net89 net119 _02191_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ net227 _04438_ _04439_ net406 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06443_ _02062_ _02076_ _02092_ _02116_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06825__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09162_ net206 _04387_ _04388_ net402 net1063 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_118_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06374_ net134 net141 net171 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_12_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08113_ net763 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[3\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__mux2_1
X_05325_ net188 _01027_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__or2_1
X_09093_ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10994__634 vssd1 vssd1 vccd1 vccd1 _10994__634/HI net634 sky130_fd_sc_hd__conb_1
X_08044_ _03575_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ net454 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05256_ _00669_ _00967_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06841__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05187_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] _00843_ _00898_
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1 vssd1 vccd1 vccd1
+ _00900_ sky130_fd_sc_hd__a22o_1
XANTENNA__07656__B _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09995_ clknet_leaf_32_wb_clk_i _00034_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_08946_ _00709_ _00710_ _04234_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared
+ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a31o_1
XANTENNA__06791__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__B2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ net435 _01389_ _02930_ _04201_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a211o_1
X_07828_ _01057_ net216 net198 _01094_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07759_ _01078_ _01513_ _01516_ _03313_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ clknet_leaf_66_wb_clk_i _00591_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09429_ _00810_ _02961_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07559__B1 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10204_ clknet_leaf_80_wb_clk_i _00208_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05367__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ clknet_leaf_57_wb_clk_i team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect
+ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.defusedGen.defusedPixel
+ sky130_fd_sc_hd__dfrtp_1
X_10066_ clknet_leaf_47_wb_clk_i _00124_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07731__B1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10968_ net608 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_31_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ net564 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978__618 vssd1 vssd1 vccd1 vccd1 _10978__618/HI net618 sky130_fd_sc_hd__conb_1
XFILLER_0_109_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05110_ net994 _00824_ _00825_ net991 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06090_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] _01772_ vssd1
+ vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold206 _00466_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold217 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[14\]
+ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold228 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[6\]
+ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05041_ _00771_ _00772_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold239 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08800_ net893 _04154_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06222__B1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] _04798_ _04803_
+ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] _02652_
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07492__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
X_05943_ net88 _01636_ _01635_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08662_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ _00707_ _04051_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__o22a_1
X_05874_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] net146
+ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__nand2_1
XANTENNA__06525__A1 _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07613_ _01647_ net102 _02762_ net147 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_89_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08593_ _03620_ _04030_ net140 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout166_A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07544_ _01646_ net102 _03101_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07475_ net951 _00824_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ net227 net405 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06426_ _02058_ _02091_ _02099_ _01693_ _02098_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06274__C net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ net206 net401 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout121_X net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06357_ net269 _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__or2_4
XFILLER_0_115_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05308_ _00993_ _00994_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__nand2_4
X_06288_ _00681_ net135 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__nor2_1
X_09076_ net208 net400 net1176 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08027_ _03564_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net389 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__mux2_1
X_05239_ _00935_ _00931_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09978_ clknet_leaf_79_wb_clk_i _00083_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_18_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] net782 net236
+ vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__mux2_1
XANTENNA__07713__B1 _03268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06449__C _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10822_ net497 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_28_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10753_ clknet_leaf_62_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\]
+ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ clknet_leaf_26_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[16\]
+ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07577__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07525__C_N net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10118_ clknet_leaf_45_wb_clk_i _00156_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10049_ clknet_leaf_63_wb_clk_i _00107_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_69_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05590_ net415 _00676_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__or3_2
XFILLER_0_19_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07104__X _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07260_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05710__D _01421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06211_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__inv_2
X_07191_ _02834_ _02838_ _02839_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07487__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06142_ net113 _01801_ _01803_ net91 _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_42_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06443__B1 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06073_ team_07_WB.instance_to_wrap.team_07.maze_clear_edge_detector.inter _00803_
+ _00804_ _00806_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__or4_2
XFILLER_0_123_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09901_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] _01777_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\] vssd1 vssd1 vccd1
+ vccd1 _04888_ sky130_fd_sc_hd__o21ai_1
X_05024_ net273 _00750_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09932__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\] _04840_ vssd1
+ vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__nand2_1
X_09763_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__inv_2
X_06975_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _02641_
+ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout283_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__nand2_1
X_05926_ net283 net280 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__or2_2
X_09694_ _04731_ _04741_ _04743_ _04730_ net1054 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a32o_1
X_08645_ _04060_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05857_ _01524_ _01533_ _01549_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout169_X net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08576_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ _03617_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_25_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05788_ _00709_ net414 _01436_ _01434_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07527_ net102 _02263_ _01708_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07458_ net451 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06409_ _01687_ _01695_ _02082_ _01647_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07389_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\] vssd1 vssd1 vccd1
+ vccd1 _02987_ sky130_fd_sc_hd__and3_1
X_09128_ net1157 net402 net209 _04362_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09059_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05788__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11021_ net388 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07844__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07336__S _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08956__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input11_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05932__X _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07162__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06476__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10805_ clknet_leaf_70_wb_clk_i _00626_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05811__C net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ clknet_leaf_57_wb_clk_i _00566_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05476__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ clknet_leaf_39_wb_clk_i _00522_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_11_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07217__A2 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ clknet_leaf_34_wb_clk_i _00462_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07754__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__B2 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__X _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06760_ _02426_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__nand2_1
XANTENNA__08866__A _00685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07770__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05711_ net481 _01423_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_125_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06691_ _02079_ _02362_ _02363_ _02210_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08430_ _03756_ _03898_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__xor2_1
X_05642_ _01348_ _01353_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_19_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08361_ _00730_ _03836_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__nand2_1
X_05573_ _01284_ _01285_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07312_ net688 net714 net731 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[2\]
+ sky130_fd_sc_hd__nor3b_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08292_ _03720_ net412 _03671_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__or3b_1
X_07243_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ _00719_ _02892_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06833__B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07174_ _02824_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07759__A3 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06125_ _01805_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06056_ net106 net141 _01645_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout302 net304 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05007_ _00738_ _00739_ _00740_ _00743_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__or4_1
Xfanout313 net315 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_2
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_2
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_4
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input3_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _04827_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__nor2_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
Xfanout368 net369 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_4
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00763_ _00780_
+ _04777_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__and4_1
X_06958_ _01691_ _02628_ _02626_ _02520_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a211o_1
XANTENNA__05068__D_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05909_ _01583_ net121 _01602_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09677_ _04731_ _04730_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
X_06889_ _02548_ _02551_ _02558_ _02559_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__and4b_1
XFILLER_0_16_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ _04047_ _04050_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__o221a_1
XANTENNA__07695__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06296__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10323__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08559_ _03650_ _03961_ _04009_ vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10521_ clknet_leaf_13_wb_clk_i _00389_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06655__B1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06743__B net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ clknet_leaf_24_wb_clk_i _00336_ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10383_ clknet_leaf_3_wb_clk_i net711 net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06958__A1 _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ net386 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07590__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07135__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05381__Y _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07686__A2 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06894__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09982__SET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10719_ clknet_leaf_56_wb_clk_i _00550_ net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07749__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06949__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07071__B1 _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06413__A3 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07930_ _03446_ _03482_ _03483_ net216 _01067_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__o32a_1
XFILLER_0_20_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07861_ net284 _03281_ _03292_ _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__or4_2
XANTENNA__05716__C _01423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09600_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] _04665_ _04675_
+ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and3_1
X_06812_ _02479_ _02481_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ net296 net119 vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__xnor2_1
XANTENNA__05385__B1 _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09531_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _04640_
+ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__nand2_1
X_06743_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ net425 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__nand2_1
XANTENNA__07126__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06828__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ net874 net202 _04604_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__o21a_1
XANTENNA__07677__A2 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06674_ _00755_ _01582_ net115 net108 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__o31a_1
X_08413_ _03753_ _03887_ _03751_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__or3b_1
X_05625_ net415 net439 _01323_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__a21o_1
X_09393_ net413 _01416_ _01477_ _04552_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10843__518 vssd1 vssd1 vccd1 vccd1 _10843__518/HI net518 sky130_fd_sc_hd__conb_1
X_08344_ net466 _03641_ _03660_ _03761_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__o31a_1
X_05556_ _01254_ _01268_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06844__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08275_ _03750_ _03753_ _03752_ _03716_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__or4b_1
XFILLER_0_117_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05487_ _00688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01199_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__o21ai_1
X_07226_ net169 _01744_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06652__A3 _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07157_ _02138_ net81 _02750_ _02807_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout201_X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06108_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__or4b_1
XFILLER_0_125_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07088_ _02134_ net82 _02732_ _02741_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a22o_1
X_06039_ net170 _01715_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__nor2_1
Xfanout110 net111 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05907__B _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_8
Xfanout132 _01577_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_6
Xfanout143 _01649_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_4
Xfanout154 net157 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_8
Xfanout165 _01719_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06168__A2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 net177 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_4
Xfanout187 _01531_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_4
Xfanout198 _01517_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_8
X_10930__579 vssd1 vssd1 vccd1 vccd1 _10930__579/HI net579 sky130_fd_sc_hd__conb_1
XFILLER_0_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09729_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\] _04767_ _04766_
+ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_83_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08937__C _01762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06738__B net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__A2 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06754__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07569__B _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10504_ clknet_leaf_27_wb_clk_i _00372_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10898__563 vssd1 vssd1 vccd1 vccd1 _10898__563/HI net563 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_59_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ clknet_leaf_44_wb_clk_i _00319_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07053__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10366_ clknet_leaf_5_wb_clk_i net749 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10297_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[10\]
+ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10245__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08856__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07659__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10946__586 vssd1 vssd1 vccd1 vccd1 _10946__586/HI net586 sky130_fd_sc_hd__conb_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05410_ _01006_ _01012_ _01026_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__nor3_1
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06390_ _02053_ _02063_ _02031_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05341_ _01028_ _01034_ _01052_ _01050_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__o31a_1
XANTENNA__07479__B _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ _03027_ _03583_ _03584_ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05272_ net421 net424 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07011_ _02656_ _02669_ _02655_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07495__A _00685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07595__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08962_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] net808
+ net445 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07913_ net105 _03381_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__o21a_1
X_08893_ _00708_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ net479 vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__o21a_1
XANTENNA__07347__A1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ _01076_ net108 vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__nand2_1
X_07775_ net431 net116 vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nand2_1
X_04987_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout363_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ net906 net205 _04634_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__o21a_1
X_06726_ _02107_ _02154_ _02260_ _02398_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05462__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08847__A1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ net956 net203 _04592_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__o21a_1
X_06657_ _02066_ _02329_ _02327_ _02328_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05608_ net440 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1
+ vccd1 vccd1 _01321_ sky130_fd_sc_hd__nor2_1
X_09376_ _04541_ net224 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__and2b_1
X_06588_ net251 _02021_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08327_ net4 _00660_ _03743_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ _00721_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__o311a_2
XFILLER_0_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05539_ _01243_ _01250_ _01251_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_90_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06724__D _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ net457 _03735_ _03736_ _03695_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07209_ _02858_ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08189_ net465 net468 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] vssd1 vssd1
+ vccd1 vccd1 _03668_ sky130_fd_sc_hd__a211o_1
X_10220_ clknet_leaf_80_wb_clk_i _00224_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05477__X _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05918__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07586__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ clknet_leaf_16_wb_clk_i net721 net322 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_7_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ clknet_leaf_67_wb_clk_i _00140_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06010__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ net624 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865__540 vssd1 vssd1 vccd1 vccd1 _10865__540/HI net540 sky130_fd_sc_hd__conb_1
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08066__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07813__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10418_ clknet_leaf_18_wb_clk_i _00309_ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_74_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08204__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10349_ clknet_leaf_33_wb_clk_i _00289_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07041__A3 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_04910_ net716 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[0\]
+ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05890_ _00716_ _01569_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nor2_1
XANTENNA__06659__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__X _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06552__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07560_ _03117_ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__or2_2
X_11009__638 vssd1 vssd1 vccd1 vccd1 _11009__638/HI net638 sky130_fd_sc_hd__conb_1
XANTENNA__05850__X _01544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06511_ _01708_ _01812_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07491_ _03045_ _03047_ _03051_ _03041_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.buttonDetect
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_61_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09230_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04435_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__nand2_1
X_06442_ _02054_ _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04907__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09161_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04384_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06373_ net200 _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__nand2_2
XFILLER_0_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08112_ net766 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05324_ net188 _01027_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__nor2_1
X_09092_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04333_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08043_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ net450 vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__mux2_1
X_05255_ net433 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05186_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] _00840_ _00898_
+ _00833_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__a22o_1
XANTENNA__07656__C _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06592__A_N _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09994_ clknet_leaf_31_wb_clk_i _00033_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10167__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07953__A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ net977 _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout199_X net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ net442 net438 vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09190__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ _01095_ net187 vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nor2_1
XANTENNA__06288__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10849__524 vssd1 vssd1 vccd1 vccd1 _10849__524/HI net524 sky130_fd_sc_hd__conb_1
X_07758_ _01066_ net214 vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06709_ _02134_ _02149_ _02375_ _02139_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07689_ _03203_ _03221_ _03246_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect
+ sky130_fd_sc_hd__or3_2
XFILLER_0_94_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09428_ _04568_ _04569_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09359_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04525_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a21o_1
XANTENNA__08048__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07559__A1 _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ clknet_leaf_83_wb_clk_i _00207_ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input41_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ clknet_leaf_43_wb_clk_i net752 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06782__A2 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ clknet_leaf_47_wb_clk_i _00123_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__07731__A1 _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06198__B _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967_ net607 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_67_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10898_ net563 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07757__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold207 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold218 _00474_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _00095_ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06470__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05040_ _00768_ _00769_ _00770_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__nand3_2
XFILLER_0_106_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06470__B2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06222__A1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ _02653_ _02654_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__nand2_1
XANTENNA__07970__A1 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__A2 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ net1148 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ net231 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
XANTENNA__07970__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07492__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05942_ _00755_ _01621_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__nor2_4
XANTENNA__05293__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ _04085_ _04087_ _04088_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a22oi_2
X_05873_ _01562_ _01564_ _01560_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a21o_1
XANTENNA__07183__C1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ _03118_ _03153_ _03169_ _02229_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__o211a_1
X_08592_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ _03618_ net871 vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07543_ net126 _01701_ net163 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10961__601 vssd1 vssd1 vccd1 vccd1 _10961__601/HI net601 sky130_fd_sc_hd__conb_1
XANTENNA__06395__Y _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout159_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07474_ net475 net1170 vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09213_ net403 _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06425_ net200 _01745_ _01663_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout326_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09144_ net325 _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06356_ net275 net278 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__nand2_4
XFILLER_0_45_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05307_ net190 _01014_ _01019_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__or3_2
XFILLER_0_44_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09075_ net323 _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__and2_1
X_06287_ _00681_ net135 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ net409 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ net291 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ _03563_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a221o_1
X_05238_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ _00948_ _00949_ _00950_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__a311o_1
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05169_ _00866_ _00880_ _00881_ _00857_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ clknet_leaf_73_wb_clk_i _00082_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__A1 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__B2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05915__B net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] net714 net236
+ vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08859_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ net295 net292 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ _04190_ vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_58_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10821_ net496 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__05931__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10752_ clknet_leaf_63_wb_clk_i _00582_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10683_ clknet_leaf_26_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[15\]
+ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07858__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05378__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06204__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10117_ clknet_leaf_45_wb_clk_i _00155_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05825__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10048_ clknet_leaf_46_wb_clk_i _00040_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataDc vssd1 vssd1 vccd1
+ vccd1 net759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06210_ net109 _01801_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06691__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__A _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07190_ _02840_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06141_ net113 _01801_ _01821_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06391__B _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06072_ net241 _01749_ _01758_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__or3_2
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ net1098 net152 net150 _04887_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a22o_1
X_05023_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net279
+ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09831_ _04840_ _04841_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\]
+ net243 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__04920__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06974_ _02641_ _02642_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__nor2_1
X_09762_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ _04785_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__and3_1
X_05925_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nand2_2
X_08713_ _04129_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ _04128_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__mux2_1
X_09693_ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08644_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nand2_1
X_05856_ _01533_ _01549_ _01524_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_68_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ _03997_ _04020_ _03996_ vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_25_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05787_ net488 _01435_ _01484_ _01433_ net490 vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07526_ _01708_ net102 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07457_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ net391 net293 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ _03029_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[6\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06408_ net124 _01701_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_40_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07388_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\] vssd1 vssd1 vccd1
+ vccd1 _02986_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_40_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09127_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06339_ net186 _01741_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__nand2_2
X_09058_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08009_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout91_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ net386 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05926__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09136__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__C1 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__B net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__B1 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08448__S net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06757__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07162__A2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ clknet_leaf_67_wb_clk_i _00625_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ clknet_leaf_57_wb_clk_i _00565_ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07588__A _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10666_ clknet_leaf_39_wb_clk_i _00521_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ clknet_leaf_35_wb_clk_i _00461_ net375 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06425__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XANTENNA__06728__A2 _02149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08866__B _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05710_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] _01417_
+ _01421_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__or4_4
XANTENNA__07770__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06690_ net88 _02148_ net249 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_125_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06667__A _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05641_ _01348_ _01353_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__or2_1
XANTENNA__06361__B1 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08360_ _01260_ _03724_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o21ai_1
X_05572_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] vssd1 vssd1 vccd1
+ vccd1 _01285_ sky130_fd_sc_hd__or3b_1
XFILLER_0_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07311_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02931_ _02934_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[2\]
+ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_3_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08291_ _03759_ _03764_ _03768_ _03630_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10622__RESET_B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06664__A1 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07173_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\] net297 _02673_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\]
+ _02823_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06416__A1 _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06124_ net117 _01797_ _01804_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06055_ net196 net201 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05006_ net32 net31 _00741_ _00742_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__or4_2
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_4
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_4
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_2
Xfanout347 net350 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_2
X_09814_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ _04826_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__and3_1
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09745_ net1036 _04776_ _04778_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout181_X net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ _02497_ _02627_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__B _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05908_ _01569_ _01578_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__xnor2_1
X_09676_ _00762_ _04710_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__nor2_2
X_06888_ net92 _02544_ _02554_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05481__A _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05839_ _01527_ _01530_ _00714_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a21oi_2
X_08627_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _04049_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08558_ _03613_ _04008_ net139 vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07509_ net166 _01739_ _02041_ _02085_ _01690_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08489_ net54 _02670_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10363__RESET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10520_ clknet_leaf_12_wb_clk_i _00388_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10451_ clknet_leaf_50_wb_clk_i _00335_ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10900__565 vssd1 vssd1 vccd1 vccd1 _10900__565/HI net565 sky130_fd_sc_hd__conb_1
XFILLER_0_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10382_ clknet_leaf_4_wb_clk_i net670 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05359__C _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05927__Y _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout94_X net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold390 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] vssd1 vssd1
+ vccd1 vccd1 net1059 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net637 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_88_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09562__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__B _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10718_ clknet_leaf_61_wb_clk_i _00549_ net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08207__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[6\]
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10245__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07860_ _03330_ _03331_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06811_ net282 _00695_ _02481_ _02480_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a31o_1
X_07791_ _03341_ _03342_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06742_ _02413_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__inv_2
X_09530_ net955 net205 _04644_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__o21a_1
XANTENNA__06397__A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__A2 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ net265 _04603_ net287 net217 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a221o_1
X_06673_ _02129_ _02312_ _02329_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__or3b_1
XANTENNA__07677__A3 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ _00048_ _03878_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a21oi_1
X_05624_ net441 _01336_ _01333_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09392_ _01415_ _01476_ net481 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10882__557 vssd1 vssd1 vccd1 vccd1 _10882__557/HI net557 sky130_fd_sc_hd__conb_1
X_08343_ net467 _03816_ _03819_ _03664_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10772__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05555_ _01266_ _01267_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout141_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout239_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08274_ net54 _00702_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__nor2_4
X_05486_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ _00689_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07225_ _02860_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07156_ _02062_ _02186_ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06107_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\] _01787_
+ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07087_ _01618_ _02214_ _02735_ _02107_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a22o_2
XFILLER_0_100_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06038_ _01668_ _01716_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout100 _01600_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout111 net112 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_2
Xfanout122 _01595_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_8
Xfanout133 net136 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_8
XFILLER_0_22_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout144 _01566_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_8
Xfanout155 net156 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_4
Xfanout166 net167 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
XANTENNA__06168__A3 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 _01544_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
X_10817__492 vssd1 vssd1 vccd1 vccd1 _10817__492/HI net492 sky130_fd_sc_hd__conb_1
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ _03455_ _03542_ _03543_ _03466_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09728_ _00772_ _00779_ _00783_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_83_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09659_ _04719_ _04718_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06876__A1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08078__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10503_ clknet_leaf_15_wb_clk_i _00371_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09578__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10434_ clknet_leaf_54_wb_clk_i _00318_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09557__S net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07053__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10365_ clknet_leaf_4_wb_clk_i net681 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05386__A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10296_ clknet_leaf_50_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[9\]
+ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05392__Y _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07106__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10285__RESET_B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06367__D net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06945__A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05340_ _01052_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05271_ net421 net422 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__xor2_2
XFILLER_0_109_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07010_ _02656_ _02669_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06680__A _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08961_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] net829
+ net444 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ net146 _03405_ _03464_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a21oi_1
X_08892_ _04211_ net952 _04209_ vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
XANTENNA__07347__A2 _00711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ _03345_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__nand2_1
X_07774_ net105 _03321_ _03326_ net106 vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__o2bb2a_1
X_04986_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
X_09513_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ net267 net289 net221 vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a211o_1
X_06725_ _02031_ _02264_ _02397_ _02128_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08847__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06656_ _02269_ _02284_ _02286_ _02265_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__o22ai_4
X_09444_ net288 _04590_ net265 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ net217 vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05607_ net442 _01314_ _01315_ _01319_ net441 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__o32a_1
XFILLER_0_47_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09375_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04538_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__and2_1
X_06587_ net250 _02021_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07022__Y _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ _03674_ _03802_ _03713_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__o21a_1
X_05538_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ _01108_ _00797_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08257_ _01296_ _01302_ net457 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a21bo_1
X_05469_ _01042_ _01051_ _01180_ _01181_ _01032_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07208_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00829_ _00943_ _02857_
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06590__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__nor2_2
XFILLER_0_104_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07139_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] net299 net394 _02790_
+ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__a22o_1
XANTENNA__05918__B net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07586__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10150_ clknet_leaf_18_wb_clk_i net713 net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05637__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ clknet_leaf_46_wb_clk_i _00139_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05482__C_N _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10983_ net623 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906__571 vssd1 vssd1 vccd1 vccd1 _10906__571/HI net571 sky130_fd_sc_hd__conb_1
XFILLER_0_92_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10417_ clknet_leaf_18_wb_clk_i _00308_ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_74_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10348_ clknet_leaf_34_wb_clk_i _00288_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06005__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__B1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10279_ clknet_leaf_81_wb_clk_i _00271_ net301 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10466__RESET_B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06510_ _02135_ _02178_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__nor2_1
X_07490_ _02034_ _02035_ _02231_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a31o_1
XANTENNA__06675__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06441_ _01734_ net164 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05512__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09160_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04384_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06372_ _01642_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08111_ net838 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[1\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05323_ _01008_ _01013_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__nor2_2
XFILLER_0_127_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09091_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04333_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ _03574_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net389 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__mux2_1
X_05254_ net433 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__04923__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05297__Y _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05185_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout104_A _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ clknet_leaf_35_wb_clk_i _00032_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ net977 _04237_ net489 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08875_ net435 _01389_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07826_ net161 _03367_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10136__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04969_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\] vssd1
+ vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
X_07757_ _01077_ net183 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06708_ net85 _02214_ _02375_ net261 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07688_ _03233_ _03237_ _03240_ _03245_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__or4_1
XANTENNA__06585__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09427_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__and2_1
X_06639_ _01596_ _01599_ _01603_ net115 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__or4_4
XFILLER_0_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09358_ net223 _04527_ _04528_ net395 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06059__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] _03683_ vssd1
+ vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09289_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04475_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_43_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05929__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08024__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ clknet_leaf_80_wb_clk_i _00206_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06767__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ clknet_leaf_43_wb_clk_i _00171_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05935__Y _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09705__B1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input34_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ clknet_leaf_47_wb_clk_i _00122_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05990__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05383__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ net606 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XANTENNA__06495__A _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10897_ net653 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_31_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07103__B net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold208 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\] vssd1 vssd1
+ vccd1 vccd1 net877 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold219 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06470__A2 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06006__Y _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06222__A2 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06990_ _01485_ _02651_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__nand2b_1
X_10915__659 vssd1 vssd1 vccd1 vccd1 net659 _10915__659/LO sky130_fd_sc_hd__conb_1
X_05941_ net96 net93 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__nand2_4
XANTENNA__07492__C _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06389__B _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05872_ _01560_ _01565_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08660_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _04047_ _04050_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ _04086_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__o221a_1
XFILLER_0_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07183__B1 _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ net144 net135 _01669_ _01672_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10363__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08591_ _03607_ _04029_ net140 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ net179 _02048_ _02887_ _01798_ _02743_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__o221a_1
XANTENNA__04918__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07473_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09212_ _04423_ _04424_ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06424_ _02043_ _02096_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ _04372_ _04373_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__and3_1
X_06355_ _02008_ _02029_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06446__C1 _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05306_ _00993_ _00994_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__or2_2
X_09074_ _04321_ _04322_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__and3_1
X_06286_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\] team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\] vssd1 vssd1 vccd1 vccd1
+ _01962_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05237_ _00907_ _00911_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ _00686_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_13_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08025_ net452 net448 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout107_X net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05168_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\]
+ _00856_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__a32o_1
XANTENNA__06749__B1 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05099_ net475 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ _00821_ _00817_ net1017 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a32o_1
X_09976_ clknet_leaf_82_wb_clk_i _00081_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08927_ net1078 net258 _04233_ vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__a21o_1
X_08858_ _03024_ net390 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07809_ net269 _03354_ _03363_ net272 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__o22a_1
XANTENNA__06586__Y _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] _04139_ net967
+ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__o21ai_1
X_10820_ net495 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_95_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10751_ clknet_leaf_64_wb_clk_i _00581_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_97_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10682_ clknet_leaf_25_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[14\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07577__C net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05378__B _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_1_0_wb_clk_i_X clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10116_ clknet_leaf_45_wb_clk_i _00154_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10386__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10047_ clknet_leaf_63_wb_clk_i net804 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 _00118_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10984__624 vssd1 vssd1 vccd1 vccd1 _10984__624/HI net624 sky130_fd_sc_hd__conb_1
XFILLER_0_86_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07114__A _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ net589 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__A_N net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07768__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06140_ _01806_ _01820_ _01807_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06071_ _01197_ _01240_ _01755_ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__or4_1
XFILLER_0_111_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05022_ net272 _00755_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07784__A _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09830_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] _04838_ net264
+ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o21ai_1
XANTENNA__05403__B1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] _04788_ _04789_
+ net244 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06973_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] net260
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] vssd1 vssd1
+ vccd1 vccd1 _02642_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08712_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ net242 vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nor2_1
X_05924_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__and2_4
X_09692_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] _04736_ vssd1 vssd1
+ vccd1 vccd1 _04742_ sky130_fd_sc_hd__and4_1
X_08643_ _01465_ _01475_ net478 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__o21a_1
X_05855_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] net180
+ net176 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] vssd1
+ vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout171_A _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout269_A net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08574_ _03617_ _04019_ net140 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__a21oi_1
X_05786_ net486 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ net474 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__o41a_1
XFILLER_0_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07525_ net159 _01689_ net165 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__or3b_1
XFILLER_0_53_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07456_ net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06407_ net126 _01702_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__nor2_2
XFILLER_0_107_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07387_ net943 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\] _02985_
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[1\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08959__A1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ net209 _04360_ _04361_ net402 net1155 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__a32o_1
X_06338_ net182 _01742_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__nor2_4
XFILLER_0_115_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09057_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__inv_2
XANTENNA__07631__A1 _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06269_ _00684_ net130 _01928_ net155 _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__o221a_1
X_08008_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09959_ clknet_leaf_79_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[28\]
+ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_95_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10968__608 vssd1 vssd1 vccd1 vccd1 _10968__608/HI net608 sky130_fd_sc_hd__conb_1
XANTENNA__07147__B1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05942__A _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__B2 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05006__X _00743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10803_ clknet_leaf_67_wb_clk_i _00624_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10734_ clknet_leaf_58_wb_clk_i _00564_ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06122__A1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10068__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ clknet_leaf_40_wb_clk_i _00520_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05389__A _00966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ clknet_leaf_35_wb_clk_i _00460_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XANTENNA__07386__B1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06667__B _02312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05640_ _01350_ _01351_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06361__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05571_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01284_ sky130_fd_sc_hd__or3b_2
XFILLER_0_129_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07310_ _02934_ _02935_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08290_ net472 net470 _03631_ _03659_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o32a_1
XANTENNA__06113__A1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07241_ _02871_ _02886_ _02891_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[3\]
+ sky130_fd_sc_hd__or3_1
XANTENNA__07498__B _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07172_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] net299 net298 team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06123_ net126 _01701_ net171 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a21o_2
XFILLER_0_124_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06416__A2 _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07613__B2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06054_ net194 net200 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__nor2_2
XFILLER_0_83_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05005_ net28 net29 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout304 net308 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_2
Xfanout315 net327 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
Xfanout326 net327 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
X_09813_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ _04825_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 _04829_ sky130_fd_sc_hd__a31o_1
Xfanout337 net351 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_2
Xfanout348 net350 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_4
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_2
XFILLER_0_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09744_ _00652_ _04777_ net244 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_20_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06956_ _02520_ _02619_ _02620_ _02622_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__or4b_1
XANTENNA__06858__A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05907_ _01590_ _01598_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__nand2_1
X_09675_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _01766_ _04709_
+ _04704_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a31o_2
XANTENNA__08877__B1 _02930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout174_X net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ _02552_ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__nor2_1
XANTENNA__05481__B _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _01249_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__and2_1
X_05838_ _01527_ _01530_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__nand2_4
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08557_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ _03612_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nand2_1
X_05769_ _01467_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\]
+ _01462_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07508_ _02036_ _02262_ net162 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06593__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08488_ net789 _03653_ _03958_ net54 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06655__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07439_ _03018_ _02984_ _03017_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[20\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_130_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07852__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ clknet_leaf_50_wb_clk_i _00334_ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09109_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04347_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ clknet_leaf_3_wb_clk_i net739 net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05937__A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold380 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_left vssd1
+ vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold391 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout87_X net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ net387 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09144__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_103_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10717_ clknet_leaf_61_wb_clk_i _00548_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10648_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[5\]
+ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09045__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06008__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10579_ clknet_leaf_60_wb_clk_i _00014_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06810_ net279 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1
+ vccd1 vccd1 _02481_ sky130_fd_sc_hd__or2_1
X_07790_ _03341_ _03342_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__nor4_1
XANTENNA__06582__B2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06741_ _02411_ _02412_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__or2_2
XANTENNA__06397__B _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__A3 _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ _04585_ _04589_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__or3_1
X_06672_ _02342_ _02344_ _02327_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a21o_1
X_08411_ net490 net462 _03715_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__o22a_1
XFILLER_0_87_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05623_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] _01316_
+ _01334_ _01335_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__a211o_1
X_09391_ net413 _01416_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08342_ net467 _03766_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__nand2_1
X_05554_ _01255_ _01265_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06637__A2 _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ _00048_ _03751_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nor2_1
X_05485_ _00688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ _00689_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07834__B2 _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout134_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ _02033_ _02758_ _02872_ _02874_ _02761_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07155_ _02134_ net81 _02741_ _02807_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout301_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07598__B1 _03144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06106_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\] _01787_
+ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__nor2_1
X_07086_ _01646_ net104 _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06037_ net974 _01633_ _01641_ _01727_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\]
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout101 _01600_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout112 _01614_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_35_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout134 net136 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_4
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout145 _03626_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_4
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout167 _01707_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
Xfanout178 _01643_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06573__A1 _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ _03376_ _03451_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nand2_1
XANTENNA__06588__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout189 _01003_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net244 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\] vssd1
+ vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and2b_1
X_06939_ _02607_ _02609_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] _04713_ _04714_
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08609_ _01202_ _04040_ _04039_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06876__A2 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _04669_ _04670_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09275__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ clknet_leaf_14_wb_clk_i _00370_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08742__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10433_ clknet_leaf_21_wb_clk_i _00317_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07053__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10364_ clknet_leaf_4_wb_clk_i net677 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10295_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[8\]
+ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09750__A1 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06498__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07106__B _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07513__B1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05270_ net422 net424 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__nand2_2
XFILLER_0_119_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07776__B net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08224__Y _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08960_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] net810
+ net444 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XANTENNA__05296__B _01008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ _03376_ _03465_ _03464_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__a21o_1
XANTENNA__07792__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ net479 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\] vssd1
+ vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09741__A1 _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07347__A3 _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ _03395_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nor2_1
XANTENNA__06555__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07773_ _03298_ _03302_ _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a21o_1
X_04985_ net718 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09512_ net912 net204 _04633_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__o21a_1
X_06724_ net254 _01714_ _01804_ _02013_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__and4_1
XFILLER_0_91_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06307__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__B1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ net480 _00813_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06655_ _00649_ net282 _00757_ _01625_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__o31a_1
XFILLER_0_8_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout251_A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout349_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05606_ net442 net439 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__nand2_1
XANTENNA__07303__Y _02930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ net397 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06586_ _01609_ _02148_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__nand2_4
XFILLER_0_47_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08325_ _03698_ _03782_ net484 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a21oi_1
X_05537_ _01248_ _01249_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08256_ _03677_ _03730_ _03732_ _03734_ _01382_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05468_ _01085_ _01127_ _01097_ _01055_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07207_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00831_ net297 team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a22o_1
XANTENNA__05758__Y _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _03646_ _03663_ _03665_ _03659_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__a31o_1
XANTENNA__06590__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05399_ _01055_ _01095_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__nor2_1
X_07138_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] net298 net297 team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ _02682_ _02707_ _02712_ _02718_ _02723_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.displayDetect
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__06794__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10080_ clknet_leaf_46_wb_clk_i _00138_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_X clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06589__Y _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06546__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06010__A3 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08299__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ net622 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_97_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05950__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09141__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06482__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10416_ clknet_leaf_18_wb_clk_i _00307_ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_115_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10347_ clknet_leaf_34_wb_clk_i _00287_ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06005__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833__508 vssd1 vssd1 vccd1 vccd1 _10833__508/HI net508 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_111_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ clknet_leaf_79_wb_clk_i _00270_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10762__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952__592 vssd1 vssd1 vccd1 vccd1 _10952__592/HI net592 sky130_fd_sc_hd__conb_1
XANTENNA__07117__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06021__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06440_ _02087_ _02112_ _02113_ _01711_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06371_ net186 _02044_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ net754 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__mux2_1
X_05322_ net426 _00991_ _01022_ _01033_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__a31o_1
X_09090_ net208 _04334_ _04335_ net397 net851 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08041_ net409 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ net291 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a221o_1
X_05253_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] net432 vssd1
+ vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05184_ _00894_ _00895_ _00896_ _00891_ _00887_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09992_ clknet_leaf_36_wb_clk_i _00031_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06776__B2 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ net980 _04235_ _04238_ vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__o21a_1
X_10890__646 vssd1 vssd1 vccd1 vccd1 net646 _10890__646/LO sky130_fd_sc_hd__conb_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08874_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\] _01372_ vssd1 vssd1
+ vccd1 vccd1 _04199_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06528__A1 _01705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07027__A _02677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _03366_ _03378_ _03376_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__or3b_2
X_07756_ _03308_ _03310_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__or2_1
XANTENNA__09478__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04968_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
X_06707_ net175 _01737_ _02013_ _02044_ net253 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_17_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07687_ _03242_ _03243_ _03244_ _03129_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__o31a_1
X_09426_ _04567_ _04570_ _04576_ _00705_ _04577_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_17_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06638_ _02303_ _02307_ _02310_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__and3_1
XANTENNA__06700__A1 _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10105__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09357_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06569_ _02050_ _02090_ _02079_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_23_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08308_ net417 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] _03785_ vssd1
+ vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_23_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09288_ net226 _04478_ _04479_ net396 net1077 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_43_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08239_ net474 _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05929__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10785__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ clknet_leaf_81_wb_clk_i _00205_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06767__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05945__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ clknet_leaf_43_wb_clk_i _00170_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10063_ clknet_leaf_47_wb_clk_i _00121_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08040__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__B1 _03269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05990__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05951__Y _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A3 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965_ net605 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_70_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10896_ net652 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_39_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold209 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[5\]
+ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06016__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06222__A3 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05940_ net99 net90 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06022__Y _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05871_ _01562_ _01564_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__and2_1
XANTENNA__07183__A1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07610_ _03098_ _03144_ _03165_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__o2bb2a_1
X_08590_ net812 _03606_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07613__A1_N _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ net179 _02048_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07472_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ net292 _03037_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[39\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09211_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ net3 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__and2_1
X_06423_ net166 _02036_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06692__Y _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ net5 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06354_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _02010_ _02027_
+ _02028_ _02026_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__04934__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06446__B1 _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05305_ _01007_ _01017_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09073_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ net4 vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06285_ _01611_ _01922_ _01960_ _01961_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.buttonHighlightDetect
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08024_ net451 net448 vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nor2_1
X_05236_ _00918_ _00923_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05167_ _00871_ _00878_ _00879_ _00864_ _00861_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10855__530 vssd1 vssd1 vccd1 vccd1 _10855__530/HI net530 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_90_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05098_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ _00817_ _00823_ net991 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a22o_1
X_09975_ clknet_leaf_79_wb_clk_i _00080_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08926_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ net234 _04228_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__and3_1
X_08857_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ net295 net292 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ _04189_ vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08371__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ _03355_ _03356_ _03362_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or3_2
XFILLER_0_58_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08788_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\]
+ _04139_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__or3_2
X_07739_ net284 _03292_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10750_ clknet_leaf_64_wb_clk_i _00580_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _04556_ _04564_ _02962_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__mux2_1
X_10681_ clknet_leaf_25_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[13\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_67_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05011__Y _00746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10115_ clknet_leaf_45_wb_clk_i _00153_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09434__X _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ clknet_leaf_46_wb_clk_i _00105_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05176__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold81 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi vssd1 vssd1
+ vccd1 vccd1 net761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05715__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07114__B _02282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07468__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ net588 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10879_ net554 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08226__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06428__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _02376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06070_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__or3b_1
XFILLER_0_112_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10839__514 vssd1 vssd1 vccd1 vccd1 _10839__514/HI net514 sky130_fd_sc_hd__conb_1
XFILLER_0_111_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05021_ net284 net278 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__nand2_8
XANTENNA__07784__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__B1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06600__B1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09760_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] _04785_ _00652_
+ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a21oi_1
X_06972_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\]
+ net260 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__and3_2
X_08711_ _01759_ _04040_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__nand3_2
X_05923_ _01590_ _01598_ net119 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a21oi_1
X_09691_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ _04736_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] vssd1 vssd1
+ vccd1 vccd1 _04741_ sky130_fd_sc_hd__a31o_1
X_08642_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04059_ _04068_ _04069_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a2bb2o_1
X_05854_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01534_
+ _01546_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ _03615_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o21ai_1
X_05785_ _01457_ _01481_ _01483_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ net138 _01688_ net165 vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07459__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10439__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net391 net293 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ _03028_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[3\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926__575 vssd1 vssd1 vccd1 vccd1 _10926__575/HI net575 sky130_fd_sc_hd__conb_1
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__04935__Y _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06406_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07386_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ net478 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_40_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09125_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ _04358_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06337_ net414 net213 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09056_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__and3_1
X_10896__652 vssd1 vssd1 vccd1 vccd1 net652 _10896__652/LO sky130_fd_sc_hd__conb_1
XFILLER_0_128_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06268_ net147 _01929_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08007_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__xor2_1
X_05219_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00932_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06199_ _01681_ _01873_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__nand2_2
XFILLER_0_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08302__C team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ clknet_leaf_82_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[25\]
+ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05782__X _01481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ net435 _01398_ _01403_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a31o_1
XANTENNA__07147__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09889_ _01775_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__nand2_1
XANTENNA__05942__B _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07698__A2 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10802_ clknet_leaf_67_wb_clk_i _00623_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08745__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ clknet_leaf_58_wb_clk_i _00563_ net333 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10664_ clknet_leaf_40_wb_clk_i _00519_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10595_ clknet_leaf_40_wb_clk_i _00459_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10151__SET_B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XANTENNA__06189__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10208__RESET_B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07138__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _00049_ _00045_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07125__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06361__A2 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05570_ _01282_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06113__A2 _00710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07240_ _02761_ _02878_ _02890_ _02781_ _02888_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a221o_1
XANTENNA__07498__C _03057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07055__A_N _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07171_ net446 team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\] net394 vssd1
+ vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06122_ net194 _01801_ _01802_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06053_ net215 net197 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05004_ net25 net24 net27 net26 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__or4_1
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 net308 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout316 net320 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_4
Xfanout327 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_4
X_09812_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] _04826_ _04828_
+ net243 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout338 net351 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_4
Xfanout349 net350 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_2
X_09743_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\]
+ _04772_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__and3_1
X_06955_ _02614_ _02618_ _02624_ _02625_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__o211a_1
XANTENNA__07129__A1 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout281_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05906_ _01590_ _01598_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__and2_2
X_09674_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _01766_ _04709_
+ _04704_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a31oi_1
X_06886_ net117 _02478_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__and2_1
XANTENNA__08877__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ _00707_ _04052_ _04048_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__a21oi_1
X_05837_ _01526_ _01529_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_85_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout167_X net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ net145 _04007_ _03965_ vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05768_ _01466_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] vssd1 vssd1 vccd1
+ vccd1 _01467_ sky130_fd_sc_hd__or3b_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07507_ net104 net165 _02036_ _02836_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08487_ _03630_ _03957_ _03653_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06593__B _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05699_ _00826_ _01411_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07438_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ _03014_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07369_ net482 _02963_ _02972_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ net208 _04346_ _04348_ net400 net1018 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__a32o_1
X_10380_ clknet_leaf_2_wb_clk_i net720 net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05937__B net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold370 team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\] vssd1 vssd1 vccd1
+ vccd1 net1039 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold381 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_left vssd1
+ vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold392 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net387 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05953__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_82_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10716_ clknet_leaf_61_wb_clk_i _00547_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05303__B1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[4\]
+ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06008__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10578_ clknet_leaf_57_wb_clk_i _00013_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06668__A1_N net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06024__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05909__A2 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08308__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _00674_ _00675_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06030__Y _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05790__B1 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06671_ _02009_ _02027_ _02170_ _02312_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__or4_1
X_08410_ _03718_ _03884_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor2_1
X_05622_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] net443
+ net440 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ _01417_ _01477_ _04550_ net230 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08341_ _03661_ _03815_ _03817_ net467 _03667_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05553_ _01255_ _01265_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08272_ net489 team_07_WB.instance_to_wrap.team_07.lcdOutput.playButtonPixel vssd1
+ vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05484_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ _01196_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07223_ net159 net107 _02872_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_A _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07154_ _02793_ _02798_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07598__A1 _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06105_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07085_ net143 _01664_ _01660_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06270__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06036_ net256 _01718_ _01721_ _01654_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__or4b_1
XFILLER_0_100_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06270__B2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout102 _01796_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout113 _01614_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_4
Xfanout124 _01595_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_8
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_2
Xfanout146 net148 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_8
XANTENNA_input1_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _01558_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_8
Xfanout168 _01685_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_87_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout179 net181 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_4
X_07987_ _03457_ _03540_ _03541_ _01679_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06573__A2 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06588__B _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ _00652_ _00780_ _00766_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__o21bai_1
X_06938_ _02515_ _02519_ _02520_ net428 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ net1175 _04717_ _04718_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__o21a_1
X_06869_ net270 _02486_ _02539_ _02537_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a31o_1
X_08608_ _01197_ _01240_ _04037_ _01755_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or4b_2
X_09588_ net1179 _04667_ net1082 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08539_ net145 _03960_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__or2_2
XFILLER_0_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10501_ clknet_leaf_14_wb_clk_i _00369_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05013__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05948__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ clknet_leaf_21_wb_clk_i _00316_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_59_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08235__C1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07589__A1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10363_ clknet_leaf_4_wb_clk_i net690 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05386__C _01021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[7\]
+ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05954__Y _01648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06131__X _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06498__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07513__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08710__B1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08474__C1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05492__A_N net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05827__A1 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08234__A _00711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__C1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07910_ net132 net121 _03378_ _03406_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__a31o_1
XANTENNA__07792__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08890_ _04210_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\]
+ _04209_ vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
XANTENNA__06689__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07841_ _01115_ net110 vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07347__A4 _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _01688_ _03321_ _03326_ _01679_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_75_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04984_ net739 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XANTENNA__05880__X _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ net267 net289 net221 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__a211o_1
X_06723_ _02134_ _02380_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07504__A1 _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09442_ net413 _01415_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__nand3b_1
X_06654_ _02272_ _02280_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05605_ net435 _01317_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__xor2_1
X_09373_ net224 _04537_ _04539_ net395 net1003 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__a32o_1
X_06585_ net88 _02148_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08324_ net774 net129 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__nor2_1
X_05536_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01239_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10096__D team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08255_ _01293_ _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__nor2_1
X_05467_ _01175_ _01177_ _01178_ _01179_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__and4b_1
XFILLER_0_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07206_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\]
+ net446 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08186_ net468 net472 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05398_ _01000_ net188 _01004_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__or3_1
XFILLER_0_132_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08768__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ net447 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07068_ _02710_ _02720_ _02722_ _02693_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_30_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07991__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06019_ net107 _01698_ _01708_ net199 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_7_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06546__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _04752_ _04753_ net1131 _04730_ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a2bb2o_1
X_10981_ net621 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05950__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08319__A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07223__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10734__RESET_B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06482__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07703__A2_N _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10415_ clknet_leaf_1_wb_clk_i _00306_ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05397__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10346_ clknet_leaf_35_wb_clk_i _00286_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_29_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10092__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872__547 vssd1 vssd1 vccd1 vccd1 _10872__547/HI net547 sky130_fd_sc_hd__conb_1
X_10277_ clknet_leaf_8_wb_clk_i _00269_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08931__A0 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08928__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06021__B _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06370_ net175 _01698_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05321_ net191 _01010_ _01021_ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08040_ net451 net448 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05252_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right _00963_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down vssd1
+ vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__or4b_4
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05183_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00890_ vssd1 vssd1
+ vccd1 vccd1 _00896_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09991_ clknet_leaf_33_wb_clk_i _00000_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06776__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ net489 _04237_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08873_ net434 _01399_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__or2_1
XANTENNA__06212__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07027__B _02681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07824_ _01697_ _03377_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04967_ net448 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
X_07755_ _01066_ net172 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06706_ _02128_ net83 _02235_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a21o_1
X_07686_ _02070_ _02278_ _02056_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05115__X _00828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ _00705_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__nor2_1
X_06637_ _01922_ _02259_ _02305_ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__o31a_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06013__A_N _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__nand2_1
X_06568_ _01647_ _01740_ _02132_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06882__A _01608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08307_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _01259_ vssd1
+ vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__nand2_1
X_05519_ _01225_ _01227_ _01230_ _01231_ _01204_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__o32a_2
X_09287_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06499_ _02163_ _02164_ _02169_ _02172_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08238_ team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\] vssd1 vssd1
+ vccd1 vccd1 _03717_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08169_ net54 net52 _00702_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__or3_2
XFILLER_0_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10200_ clknet_leaf_80_wb_clk_i _00204_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07964__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ clknet_leaf_43_wb_clk_i _00169_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05945__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10062_ clknet_leaf_47_wb_clk_i _00120_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08748__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05961__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10964_ net604 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__05025__X _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06152__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ net651 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07888__A _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06016__B net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07955__A1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ clknet_leaf_24_wb_clk_i net686 net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06032__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__A1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05870_ _01534_ _01563_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__xor2_1
XANTENNA__06967__A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07183__A2 _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07540_ _01618_ _01623_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__nand2_2
XFILLER_0_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07471_ _00706_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ net392 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09210_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ net3 vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nor2_1
X_06422_ net104 net166 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06694__B2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09141_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ net5 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06353_ _00709_ net270 _02009_ net120 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_20_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06446__A1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05304_ _01012_ _01016_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ net4 vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__or2_1
X_06284_ net86 _01634_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ net489 _03561_ _00796_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__mux2_1
X_05235_ _00887_ _00891_ _00892_ _00893_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10959__599 vssd1 vssd1 vccd1 vccd1 _10959__599/HI net599 sky130_fd_sc_hd__conb_1
X_05166_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06749__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__B2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05097_ net475 _00814_ _00821_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__and3_2
X_09974_ clknet_leaf_83_wb_clk_i _00079_ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07038__A _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ net861 net234 _04231_ _04232_ vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout197_X net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _03024_ net390 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08371__A1 _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _03357_ _03358_ _03360_ _03361_ _03359_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05999_ net133 net128 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__nand2_4
X_08787_ _04145_ _04146_ net192 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07044__Y _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ _03289_ _03291_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__or2_1
X_07669_ net159 _01688_ _03198_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07331__C1 _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09408_ team_07_WB.instance_to_wrap.team_07.sck_rs_enable _04563_ net411 team_07_WB.instance_to_wrap.team_07.sck_fl_enable
+ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a211o_1
XANTENNA__06685__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ clknet_leaf_25_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[12\]
+ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06117__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05021__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05956__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09387__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10114_ clknet_leaf_44_wb_clk_i _00152_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10045_ clknet_leaf_63_wb_clk_i _00104_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi
+ sky130_fd_sc_hd__dfxtp_1
Xhold60 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__A2 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05691__A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold71 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold82 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05176__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold93 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc vssd1 vssd1 vccd1
+ vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07454__A_N net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10947_ net587 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_86_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10878_ net553 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08226__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06428__A1 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10921__665 vssd1 vssd1 vccd1 vccd1 net665 _10921__665/LO sky130_fd_sc_hd__conb_1
X_10878__553 vssd1 vssd1 vccd1 vccd1 _10878__553/HI net553 sky130_fd_sc_hd__conb_1
XANTENNA_2 team_07_WB.instance_to_wrap.team_07.borderGen.synchronized_rectangle_pixel
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05020_ net275 net274 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__nor2_2
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06971_ _00716_ net260 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05872__Y _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01243_ _04035_ net242 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a31o_1
X_05922_ _01597_ _01604_ net111 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__and3_4
X_09690_ _00699_ _04739_ _04740_ net246 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a22oi_1
X_05853_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01546_
+ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__and2_1
X_08641_ net455 _04067_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05784_ _00792_ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\] _01481_
+ _01482_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__or4_1
X_08572_ _04013_ _04018_ _03996_ vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__o21a_1
X_07523_ net162 _02836_ _01678_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_25_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07454_ net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04945__A team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06405_ _00635_ net279 _00749_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__and3_4
X_07385_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\] net230 vssd1
+ vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[0\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06419__A1 _02074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09124_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ _04358_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__or2_1
XANTENNA__07616__B1 _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06336_ net414 net177 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07092__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09055_ net946 net407 net248 _04306_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__a22o_1
X_06267_ _01943_ _01940_ net251 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__and3b_1
XFILLER_0_60_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05218_ _00929_ _00930_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1 vssd1 vccd1 vccd1
+ _00931_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_13_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08006_ _03554_ _03555_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06224__X _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07694__C _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06198_ _01656_ _01829_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05149_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1 vssd1 vccd1 vccd1
+ _00862_ sky130_fd_sc_hd__mux2_1
XANTENNA__08041__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09957_ clknet_leaf_79_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[24\]
+ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_08908_ net974 _04219_ net259 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__o21a_1
X_09888_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] _01774_ vssd1
+ vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
XANTENNA__07147__A2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ net814 _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07698__A3 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05016__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ clknet_leaf_70_wb_clk_i _00622_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10732_ clknet_leaf_58_wb_clk_i _00562_ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__A _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10663_ clknet_leaf_40_wb_clk_i _00518_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10594_ clknet_leaf_35_wb_clk_i _00458_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08761__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07083__A1 _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07083__B2 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10990__630 vssd1 vssd1 vccd1 vccd1 _10990__630/HI net630 sky130_fd_sc_hd__conb_1
XFILLER_0_120_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06013__C _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10028_ _00048_ _00635_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_37_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07125__B _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10028__CLK _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07170_ _02819_ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06121_ _01800_ _01801_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05867__Y _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06052_ net210 net194 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__nor2_4
XANTENNA__06821__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05003_ net18 net17 net15 net16 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout306 net308 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_4
X_09811_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ _00657_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a21oi_1
Xfanout317 net320 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_4
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_4
X_09742_ net245 _04774_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__nor2_1
X_06954_ net211 _02510_ _02616_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07129__A2 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05905_ _01585_ _01589_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09673_ _04727_ _04728_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__nor2_1
X_06885_ _02546_ _02547_ _02549_ _02555_ _02473_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__o221a_1
XANTENNA__06888__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ net455 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__mux4_1
X_05836_ _01521_ _01528_ _01513_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_68_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07603__X _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10099__D team_07_WB.instance_to_wrap.team_07.memGen.buttonHighlightDetect
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ _03612_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nand2_1
X_05767_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] vssd1 vssd1 vccd1
+ vccd1 _01466_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07506_ _01632_ _02181_ _03063_ _03064_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_37_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08486_ net471 _03631_ _03955_ _03956_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__o211a_1
X_05698_ _01195_ _01410_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07437_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ _03013_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] vssd1
+ vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07986__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07368_ net482 _02963_ _02970_ _02973_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[1\]
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_131_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09107_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__inv_2
XANTENNA__07065__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06319_ net194 _01977_ _01979_ _01978_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a31o_1
X_07299_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ _01321_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__a31o_1
X_10974__614 vssd1 vssd1 vccd1 vccd1 _10974__614/HI net614 sky130_fd_sc_hd__conb_1
X_09038_ net248 _04293_ _04295_ net407 net1156 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] vssd1 vssd1
+ vccd1 vccd1 net1029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1040 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold382 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11000_ net386 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
Xhold393 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] vssd1 vssd1
+ vccd1 vccd1 net1062 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06576__B1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05953__B _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07226__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06130__A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10341__RESET_B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07828__B1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10715_ clknet_leaf_61_wb_clk_i _00546_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10646_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[3\]
+ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10577_ clknet_leaf_9_wb_clk_i _00445_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06024__B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06567__B1 _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06040__A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08859__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05790__B2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10082__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06670_ _02009_ _02313_ _02027_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__a21o_1
XANTENNA__06975__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10011__RESET_B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05621_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] net443
+ _00679_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08340_ _03660_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__or2_1
X_05552_ _01256_ _01264_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ _03718_ _03748_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__o21ba_1
X_05483_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07222_ _01645_ _01744_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07153_ _02802_ _02805_ _02799_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06104_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\]
+ _01786_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__or3_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ net253 net170 _02154_ _01663_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06035_ _01654_ _01719_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout103 _01796_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_35_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout114 _01614_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout125 net127 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout136 _01576_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_4
XANTENNA_fanout489_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout158 net161 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_87_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout169 _01681_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_4
X_07986_ net257 _03379_ _03387_ _03406_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_52_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ _04733_ _04764_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__nor2_1
X_06937_ _02514_ _02592_ _02515_ _02513_ _02522_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09656_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] _04717_ _04716_
+ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a21oi_1
X_06868_ _02536_ _02538_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__nor2_1
X_08607_ _00688_ _04037_ _04038_ _04039_ vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__o2bb2a_1
X_05819_ _00713_ _01501_ _01504_ _01512_ _01492_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__a2111o_4
X_09587_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ _04667_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__and3_1
X_06799_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _02467_ _02469_
+ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a21oi_2
X_08538_ net815 _03607_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08469_ net457 _01301_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10500_ clknet_leaf_14_wb_clk_i _00368_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10824__499 vssd1 vssd1 vccd1 vccd1 _10824__499/HI net499 sky130_fd_sc_hd__conb_1
X_10431_ clknet_leaf_53_wb_clk_i _00315_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05948__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08324__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10362_ clknet_leaf_5_wb_clk_i net697 net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06261__A2 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10293_ clknet_leaf_49_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[6\]
+ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout92_X net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05964__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06549__B1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06498__C _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07513__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05637__A_N net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05827__A2 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10629_ clknet_leaf_39_wb_clk_i _00493_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05874__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06689__B net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _01050_ net119 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__xnor2_1
XANTENNA__05593__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06555__A3 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _03303_ _03324_ _03325_ _03306_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04983_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
X_09510_ net894 net204 _04632_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__o21a_1
X_06722_ _02140_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07504__A2 _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _04549_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__and2_1
X_06653_ _02311_ _02325_ net420 net419 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05604_ _01315_ net442 _01314_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__or3b_1
X_09372_ _04538_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07313__B team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06584_ _01618_ _02147_ _02175_ _02257_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ net959 _03800_ net129 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05535_ _01194_ _01247_ _01245_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ net458 _01304_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05466_ _01033_ _01052_ net432 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_31_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07205_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] net298 _00942_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_43_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08185_ net468 net473 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and2_1
X_05397_ _01000_ net189 _01004_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__nor3_1
XFILLER_0_131_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07136_ _02730_ _02753_ _02755_ _02778_ _02789_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[0\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10463__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07067_ _02689_ _02709_ _02715_ _02110_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06018_ _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06546__A3 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ _01113_ net183 net169 vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__o21a_1
XANTENNA__06951__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\] _04750_ _04731_
+ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10980_ net620 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__08299__A3 _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _04702_ _00761_
+ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__o21a_1
XANTENNA__06703__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05506__B2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07223__B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05024__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06482__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ clknet_leaf_1_wb_clk_i _00305_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\]
+ sky130_fd_sc_hd__dfstp_4
XTAP_TAPCELL_ROW_115_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10703__RESET_B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10345_ clknet_leaf_35_wb_clk_i _00285_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__B1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ clknet_leaf_4_wb_clk_i _00268_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08220__D team_07_WB.instance_to_wrap.team_07.displayPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06942__B1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06021__C _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05320_ net190 _01025_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05251_ _00658_ _00794_ _00963_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__nor3_4
XANTENNA__07670__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05182_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00886_ vssd1 vssd1
+ vccd1 vccd1 _00895_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05875__Y _01569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09990_ clknet_leaf_36_wb_clk_i _00030_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08941_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ _04234_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ net439 net832 net242 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07823_ _01697_ _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__nor2_1
X_07754_ _01066_ net172 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__nand2_1
X_04966_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XANTENNA__07489__A1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06705_ _02013_ _02073_ _02370_ _02371_ _02377_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a41o_1
X_07685_ _01739_ _02036_ _03198_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout354_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _04571_ _04575_ _04576_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06636_ _02108_ _02259_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__or3b_1
XANTENNA__06161__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10458__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ net996 net395 net223 _04526_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06567_ _02051_ _02121_ _02240_ _02067_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08306_ net488 _03783_ _03713_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05518_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\] _01222_
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__mux2_1
X_09286_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__nand2_1
X_06498_ net199 net249 _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05131__X _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08237_ net462 _03714_ _03715_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05449_ _01071_ _01161_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08168_ _03630_ _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07119_ _02771_ _02772_ _02769_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_63_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08099_ net989 net229 _03595_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10130_ clknet_leaf_43_wb_clk_i _00168_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06403__A _02074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10061_ clknet_leaf_47_wb_clk_i _00119_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05019__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05961__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10963_ net603 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08209__A_N net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10894_ net650 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07888__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07652__A1 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ clknet_leaf_24_wb_clk_i net725 net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06313__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10259_ clknet_leaf_7_wb_clk_i _00251_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06032__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07470_ net1143 net292 _03036_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[38\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06421_ _02063_ _02094_ _02080_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06694__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09140_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ _04371_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06352_ net99 _01616_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_6_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_20_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05303_ _01013_ _01015_ net191 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__a21oi_1
X_09071_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ _04320_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__o2111ai_1
XANTENNA__06446__A2 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07643__A1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06283_ _01610_ net271 _01957_ _01959_ net100 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08022_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _03561_ sky130_fd_sc_hd__or2_1
X_05234_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] net299 _00830_ vssd1
+ vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__A1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05165_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07319__A _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05096_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00819_ vssd1 vssd1 vccd1
+ vccd1 _00822_ sky130_fd_sc_hd__nand2_1
X_09973_ clknet_leaf_80_wb_clk_i _00078_ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_90_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06223__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ _04228_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__and2_1
XANTENNA__07159__B1 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__X team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net391 net291 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ _04188_ vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ _01048_ net116 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08786_ net1012 _04139_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__nand2_1
X_05998_ net132 net121 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__nor2_4
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _03289_ _03291_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__nor2_1
X_04949_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07668_ _02081_ _02260_ _02277_ _01729_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06134__A1 _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06893__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07331__B1 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09407_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ _00818_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_45_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06619_ _01812_ _02283_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__or2_1
XANTENNA__06685__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ _03139_ _03141_ _03157_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09338_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07634__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10366__RESET_B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09269_ _04419_ _04429_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05021__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08613__A _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05956__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ clknet_leaf_45_wb_clk_i _00151_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08759__S net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05972__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _00064_ _00642_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold50 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_76_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07165__A3 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05691__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold72 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\] vssd1 vssd1
+ vccd1 vccd1 net741 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold83 _00172_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\] vssd1
+ vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10946_ net586 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10877_ net552 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05716__B_N _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06428__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07625__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_3 team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06600__A2 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06970_ _02570_ _02583_ _02601_ _02640_ _02572_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__05882__A _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05921_ _01583_ net121 _01613_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a21o_2
X_08640_ net455 _04067_ _04066_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__o21ai_1
X_05852_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] net176
+ _01545_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09073__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ _03616_ _04017_ net139 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a21oi_1
X_05783_ _00777_ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\] vssd1 vssd1 vccd1
+ vccd1 _01482_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07522_ _02785_ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07453_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net391 net293 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ _03025_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[2\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06404_ _02068_ _02077_ _02066_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07384_ net410 _01475_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__nor2_1
X_09123_ net209 _04357_ _04359_ net400 net981 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__a32o_1
XANTENNA__05122__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06419__A2 _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07616__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06335_ net87 _02009_ net101 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07616__B2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09054_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ _04301_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a31o_1
XANTENNA__07092__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06266_ _01924_ _01925_ _01932_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08005_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__xor2_1
X_05217_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout105_X net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06197_ _01659_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08041__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05148_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00861_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09956_ clknet_leaf_82_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[7\]
+ net300 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_05079_ _00803_ _00804_ _00806_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear
+ sky130_fd_sc_hd__nor3_1
X_08907_ _01397_ _01405_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__nor2_1
X_09887_ net844 net151 net149 _04879_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ _04178_ _04179_ _04144_ vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08769_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] net776 net239 vssd1
+ vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10800_ clknet_leaf_70_wb_clk_i _00621_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05016__B net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ clknet_leaf_58_wb_clk_i _00561_ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07855__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__B _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10662_ clknet_leaf_41_wb_clk_i _00517_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07607__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ clknet_leaf_37_wb_clk_i _00457_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05967__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08032__A1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08032__B2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XANTENNA__06043__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06013__D _01705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10027_ clknet_leaf_52_wb_clk_i _00004_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06310__B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10929_ net578 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
X_10845__520 vssd1 vssd1 vccd1 vccd1 _10845__520/HI net520 sky130_fd_sc_hd__conb_1
XFILLER_0_85_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06120_ _01668_ net102 _01798_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06051_ _01678_ net142 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__nand2_2
XANTENNA__06044__Y _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05002_ net21 net20 net23 net22 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_2
X_09810_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] net243 vssd1
+ vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__nor2_1
XANTENNA__05883__Y _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 net320 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
Xfanout329 net332 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07782__B1 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _04767_ _04774_ _04775_ net245 net1120 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__a32o_1
X_06953_ _02621_ _02622_ _02623_ _02619_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a31o_1
X_05904_ _01585_ net122 _01589_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a21o_4
X_10932__581 vssd1 vssd1 vccd1 vccd1 _10932__581/HI net581 sky130_fd_sc_hd__conb_1
X_09672_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\]
+ _04725_ _04716_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a31o_1
X_06884_ _02551_ _02552_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05117__A _00685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net455 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__nand2b_1
X_05835_ _01521_ _01528_ _01513_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_85_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06682__C_N _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ _03611_ net1114 vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__o21ai_1
X_05766_ _01461_ _01462_ _01463_ _01464_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__and4b_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07505_ _01619_ _01922_ _02217_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_18_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08485_ _03667_ _03953_ _03925_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05697_ _00687_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01252_
+ _01409_ _00962_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__o311a_1
XFILLER_0_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ net963 _03014_ _03016_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[19\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07367_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09106_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__and3_1
X_06318_ _01964_ _01971_ _01970_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07065__A2 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07298_ _02926_ _02927_ _01321_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[3\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05076__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09037_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06249_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] net456 vssd1 vssd1
+ vccd1 vccd1 _01926_ sky130_fd_sc_hd__or2_2
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold350 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 net1019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold361 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\] vssd1 vssd1 vccd1
+ vccd1 net1030 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold372 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\] vssd1
+ vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold394 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout82_A _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06411__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ net464 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06130__B _01692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05027__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10829__504 vssd1 vssd1 vccd1 vccd1 _10829__504/HI net504 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_103_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07828__B2 _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10714_ clknet_leaf_60_wb_clk_i _00545_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08772__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06500__A1 _02139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10645_ clknet_leaf_38_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[2\]
+ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05968__Y _01662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10576_ clknet_leaf_9_wb_clk_i _00444_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05984__X _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10765__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_127_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06319__A1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05790__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10469__RESET_B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__B _02641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05620_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] _01316_
+ _01332_ _00679_ _00680_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05551_ _01262_ _01263_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08270_ _00048_ _03715_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or2_1
X_05482_ _01194_ _01192_ _01190_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__or3b_2
XANTENNA__10286__Q team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07221_ _01645_ _01744_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07152_ net107 _01710_ _02767_ _02804_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06103_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ _01784_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07083_ _02065_ net82 _02732_ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06034_ _01662_ _01723_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout104 _01694_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06558__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout115 net116 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_4
Xfanout137 _01648_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 _01567_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_6
Xfanout159 net161 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_4
X_07985_ _03374_ _03539_ _03460_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09724_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\] net246 _04761_
+ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_52_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06936_ _02521_ _02592_ _02595_ _02606_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__or4_1
XANTENNA__07507__B1 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09655_ _04703_ _04710_ _04714_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06867_ net280 _02474_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout172_X net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _00688_ _01242_ _01755_ _04037_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__a31o_1
X_05818_ _00712_ _01496_ _01510_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__or3_1
X_09586_ net1087 _04667_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__xor2_1
X_06798_ _00696_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02469_ sky130_fd_sc_hd__and2_1
XANTENNA__05533__A2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07062__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ _03994_ _03993_ net1006 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05749_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] vssd1 vssd1 vccd1
+ vccd1 _01448_ sky130_fd_sc_hd__or3_2
XFILLER_0_65_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08468_ net457 _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07419_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] _03004_
+ net477 vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08399_ net485 _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10430_ clknet_leaf_54_wb_clk_i _00314_ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06406__A _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05310__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10361_ clknet_leaf_5_wb_clk_i _00038_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06261__A3 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ clknet_leaf_49_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[5\]
+ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05964__B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\] vssd1 vssd1 vccd1
+ vccd1 net860 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06412__Y _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__A _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07513__A3 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06721__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05919__A2_N _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05204__B _00846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05698__Y _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ clknet_leaf_39_wb_clk_i _00492_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10559_ clknet_leaf_13_wb_clk_i _00427_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__A1 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05874__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06689__C net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06051__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ net296 net172 vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__xnor2_1
X_04982_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
X_06721_ net174 _01702_ _02014_ _02393_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09440_ net922 net218 net287 _04588_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__a22o_1
X_06652_ _02129_ _02287_ _02312_ _02319_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__o311a_1
X_05603_ net443 _00679_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__nor2_1
X_09371_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04533_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06583_ net84 _02179_ _02206_ _02239_ _02256_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a2111o_1
X_08322_ _03753_ _03799_ _03769_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05534_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _00793_ _00794_ _01231_ _01246_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08253_ net459 _03731_ net458 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05465_ _00982_ _01074_ _01091_ _01073_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_31_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout132_A _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00829_ net394 _02854_
+ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08184_ net465 net468 _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06226__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05396_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ _01108_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07135_ _01646_ _02783_ _02784_ _02754_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06779__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ net121 _01676_ net167 _02716_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06017_ net158 net166 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_54_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06400__B1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08940__A2 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _01113_ net172 _03371_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a21o_1
X_09707_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ _04749_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and3_1
X_06919_ _02576_ _02577_ _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__o21ba_1
X_07899_ _03383_ _03386_ _03453_ _03452_ _03387_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__o32a_1
X_09638_ _00654_ _00764_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__and2_1
XANTENNA__06703__A1 _02066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__B2 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09569_ _04612_ _04626_ _04657_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06407__Y _02081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10413_ clknet_leaf_1_wb_clk_i _00304_ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05975__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10344_ clknet_leaf_56_wb_clk_i _00284_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10275_ clknet_leaf_7_wb_clk_i _00267_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08695__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08447__A1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06972__C net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05250_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__or3_2
XANTENNA__07670__A2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06046__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05181_ _00892_ _00893_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06630__B1 _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ net1041 _04234_ _04236_ vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06052__Y _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08871_ net441 net795 net242 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
X_07822_ _01095_ net154 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ _01067_ net171 vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__nor2_1
X_04965_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] vssd1
+ vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ _02271_ _02373_ _02374_ _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__and4_1
X_07684_ _03131_ _03172_ _03241_ _03126_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__o31a_1
XANTENNA__07489__A2 _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ _00808_ _04567_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nand2_1
X_06635_ _02266_ _02293_ _02300_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_59_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout347_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09354_ _04524_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06566_ net199 _02124_ _02194_ _02097_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06508__X _02182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ net484 _03776_ _03781_ _03770_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__o31a_1
X_05517_ _01204_ _01229_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__nand2_1
X_09285_ net226 _04476_ _04477_ net396 net867 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06497_ _01646_ _01734_ _01660_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08236_ net410 _03561_ net489 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05448_ _01104_ _01107_ _01100_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08870__S net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05672__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08167_ net54 net52 net53 _03627_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__o31a_1
XANTENNA__04970__Y _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05379_ _00970_ _01058_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07118_ net273 _02106_ net81 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08098_ _03601_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ _03594_ vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06621__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07049_ _01921_ _02258_ net83 net261 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10060_ clknet_leaf_46_wb_clk_i net760 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataDc
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_110_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05019__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08110__S team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10962_ net602 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XFILLER_0_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10893_ net649 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07521__Y _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06418__X _02092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07652__A2 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ clknet_leaf_25_wb_clk_i net716 net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_130_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10258_ clknet_leaf_7_wb_clk_i _00250_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10189_ clknet_leaf_74_wb_clk_i net730 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07712__X _03268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__B1 _02250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07340__A1 _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07340__B2 _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06420_ _02084_ _02093_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06351_ net257 _02017_ _02024_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06047__Y _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05302_ _00996_ _01014_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__or2_2
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09070_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04319_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__o21a_1
X_06282_ net124 _01958_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07643__A2 _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ _03560_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[1\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05233_ _00939_ _00940_ _00945_ _00834_ _00832_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__a32o_1
X_05164_ _00854_ _00875_ _00876_ _00847_ _00845_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05095_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00819_ vssd1 vssd1 vccd1
+ vccd1 _00821_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ clknet_leaf_72_wb_clk_i _00077_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07319__B _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06223__B _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06666__A1_N net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ net235 _04229_ _04231_ vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__o22a_1
XANTENNA__07159__A1 _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08854_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ net293 net389 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__a22o_1
XANTENNA__07564__D1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ _01049_ net118 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08785_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] _04139_ vssd1
+ vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__or2_1
X_05997_ net137 net168 _01688_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__and3_2
XFILLER_0_137_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ net277 _01105_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04948_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
X_07667_ _03065_ _03223_ _03224_ _03095_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__A1 _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ net960 _04562_ _04558_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06618_ _02129_ _02281_ _02287_ _02067_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__o221a_1
X_07598_ _03098_ _03143_ _03144_ _03148_ _03156_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__o221a_1
X_10862__537 vssd1 vssd1 vccd1 vccd1 _10862__537/HI net537 sky130_fd_sc_hd__conb_1
XANTENNA__10379__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09337_ net223 _04512_ _04513_ net395 net1154 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a32o_1
X_06549_ _00758_ net87 net98 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a21o_1
XANTENNA__07501__C _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ _04418_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07634__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ net412 _03697_ net487 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09199_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04378_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09387__A2 _01475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10112_ clknet_leaf_44_wb_clk_i _00150_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10043_ _00063_ _00641_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ sky130_fd_sc_hd__dfxtp_2
Xhold40 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold73 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _00113_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10945_ net585 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10876_ net551 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__06530__C1 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07873__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05884__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06308__B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05987__X _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05212__B _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07625__A2 _03079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08050__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05920_ _01583_ net121 _01613_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a21oi_4
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05882__B _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05851_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] _01536_
+ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08570_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ _03615_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__nand2_1
X_05782_ _01477_ _01479_ _01457_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__or3b_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07521_ _01655_ _01685_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07452_ net293 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06403_ _02074_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07383_ _02965_ _02983_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _04358_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__inv_2
XANTENNA__05122__B team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06334_ _00751_ _01620_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__or2_4
XANTENNA__07616__A2 _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05627__B2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ net1159 net407 net248 _04305_ vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06265_ net212 _01926_ _01930_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout212_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08004_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__xor2_1
X_05216_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06196_ net212 _01656_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05147_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] _00859_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_4
XFILLER_0_111_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09955_ clknet_leaf_80_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[6\]
+ net302 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05078_ _00672_ net429 _00696_ net425 _00805_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__a221o_1
X_08906_ _00682_ _04218_ net242 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__a21oi_1
X_09886_ _01774_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nand2_1
X_08837_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\]
+ _04142_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__or3_1
XANTENNA__07552__A1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08768_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] net787 net240 vssd1
+ vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07719_ _01065_ _01590_ _01598_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_64_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _01240_ _04064_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ clknet_leaf_58_wb_clk_i _00560_ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07512__B _03070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05313__A _01008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10661_ clknet_leaf_19_wb_clk_i _00516_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_101_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06128__B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10592_ clknet_leaf_36_wb_clk_i _00456_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07607__A2 _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05967__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05983__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06043__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11012__639 vssd1 vssd1 vccd1 vccd1 _11012__639/HI net639 sky130_fd_sc_hd__conb_1
X_10026_ clknet_leaf_48_wb_clk_i _00003_ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05207__B _00844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10949__589 vssd1 vssd1 vccd1 vccd1 _10949__589/HI net589 sky130_fd_sc_hd__conb_1
XFILLER_0_85_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10928_ net577 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09048__B2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10859_ net534 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06050_ _01679_ _01698_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__nor2_4
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06054__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05001_ _00734_ _00735_ _00736_ _00737_ vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__or4_2
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout308 net327 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_2
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07782__A1 _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] _04772_ vssd1
+ vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__or2_1
X_06952_ net160 _02504_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__or3b_1
.ends

