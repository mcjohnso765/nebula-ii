/*
* This is a template for your top level test bench!
* You are responsible for having a test bench for your top
* level design. Otherwise, your design will not be part
* of the tape-out.
*
* Please also include test benches for your team_04_WB
* and team_04_Wrapper modules, if needed to verify
* interfacing with the Wishbone Bus.
*
* The command to run this test bench is:
* make tbsim-source-team_04-team_04
*/

`timescale 1 ns / 1 ps

module team_04_tb();

    logic tb_clk, nrst; //clock and reset signals

endmodule
