* NGSPICE file created from team_10_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt team_10_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__2479__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3155_ _1564_ _1583_ _0906_ _1562_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__o2bb2a_1
X_2106_ team_10_WB.instance_to_wrap.dispFSM.guesses\[6\] net114 net140 net642 vssd1
+ vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__o22a_1
X_3086_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _1537_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[79\] sky130_fd_sc_hd__mux2_1
X_2037_ team_10_WB.instance_to_wrap.dispFSM.guesses\[75\] net112 net138 team_10_WB.instance_to_wrap.dispFSM.msg\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout162_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3443__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3988_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[25\]
+ _0056_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2939_ net213 net151 net120 net668 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[44\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4502__313 vssd1 vssd1 vccd1 vccd1 _4502__313/HI net313 sky130_fd_sc_hd__conb_1
XANTENNA__2954__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2190__A team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4108__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4609_ net383 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4258__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3924__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3425__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3911_ net290 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1987__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3842_ net272 vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2936__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3773_ net263 vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ _1351_ team_10_WB.instance_to_wrap.clock_div.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _1355_ sky130_fd_sc_hd__a31o_1
X_2655_ _1308_ _1310_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4325_ clknet_leaf_14_wb_clk_i _0715_ _0314_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[48\]
+ sky130_fd_sc_hd__dfstp_1
X_2586_ _0888_ _0902_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__nand2_1
XANTENNA__4400__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3045__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout138 net142 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
Xfanout127 net128 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
Xfanout116 _0913_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dlymetal6s2s_1
X_4256_ clknet_leaf_0_wb_clk_i _0650_ _0245_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.green
+ sky130_fd_sc_hd__dfrtp_1
X_3207_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] _1621_ vssd1 vssd1 vccd1
+ vccd1 _1622_ sky130_fd_sc_hd__and2_1
X_4187_ clknet_leaf_12_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[49\]
+ _0176_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[49\] sky130_fd_sc_hd__dfrtp_1
X_3138_ _1549_ _1567_ _1568_ _1551_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1
+ vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_107_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4647__415 vssd1 vssd1 vccd1 vccd1 _4647__415/HI net415 sky130_fd_sc_hd__conb_1
XANTENNA__3416__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2185__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3069_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__mux2_1
XANTENNA__4173__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3744__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] vssd1 vssd1 vccd1 vccd1
+ net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\] vssd1 vssd1 vccd1
+ vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] vssd1 vssd1 vccd1 vccd1
+ net637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2794__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_124_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3407__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3919__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1969__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4423__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ net500 net132 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\]
+ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3343__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2371_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] _1084_ _1144_
+ _1145_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__o22a_1
X_4110_ clknet_leaf_20_wb_clk_i net491 _0109_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_4041_ clknet_leaf_21_wb_clk_i _0526_ _0082_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_142_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1902__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_151_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3825_ net288 vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
XANTENNA__2452__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3756_ net292 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2707_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[2\] vssd1 vssd1 vccd1 vccd1 _1345_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3687_ net250 vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__inv_2
X_2638_ _0922_ _0925_ _0935_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] _0975_
+ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__o221a_1
X_2569_ net222 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] net226 vssd1
+ vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_160_Left_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4308_ clknet_leaf_21_wb_clk_i net612 _0297_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4168__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4239_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[3\]
+ _0228_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4446__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1940_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] net146 vssd1 vssd1 vccd1
+ vccd1 _0863_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1871_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] vssd1 vssd1 vccd1 vccd1
+ _0796_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4590_ net453 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_3610_ net282 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3541_ net245 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3472_ team_10_WB.instance_to_wrap.dispFSM.guesses\[79\] _1715_ _1842_ _0821_ vssd1
+ vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2423_ net462 net129 vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__or2_1
XANTENNA__3963__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2354_ _1126_ _1128_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4319__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2285_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _1063_ _1064_ _1066_ vssd1
+ vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2447__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4024_ clknet_leaf_0_wb_clk_i net524 _0071_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4469__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3559__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3808_ net262 vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3739_ net276 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3188__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3986__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3932__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2070_ team_10_WB.instance_to_wrap.dispFSM.guesses\[42\] net111 net136 net675 vssd1
+ vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3482__B1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2037__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2972_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] _0835_ net161 vssd1 vssd1 vccd1
+ vccd1 _1487_ sky130_fd_sc_hd__a41o_1
XFILLER_0_173_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1923_ net4 net5 net299 vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_192_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4642_ net410 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ net448 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3524_ net232 vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_151_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3455_ team_10_WB.instance_to_wrap.host_row2\[54\] net171 net168 team_10_WB.instance_to_wrap.host_row2\[78\]
+ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload27_A clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4141__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2406_ team_10_WB.instance_to_wrap.clock_div.count\[19\] team_10_WB.instance_to_wrap.clock_div.count\[18\]
+ team_10_WB.instance_to_wrap.clock_div.count\[21\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__or4_1
X_3386_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] net169 _1727_ team_10_WB.instance_to_wrap.dispFSM.guesses\[43\]
+ _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_110_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2337_ _0809_ _0866_ _1093_ _0811_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__a22oi_1
X_2268_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0800_ net214 _0792_ vssd1
+ vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_162_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4291__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4007_ clknet_leaf_26_wb_clk_i _0495_ net239 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2199_ _0984_ _0987_ _0975_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2640__B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold41 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] vssd1 vssd1 vccd1 vccd1
+ net497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 team_10_WB.instance_to_wrap.message_reg.msg\[4\] vssd1 vssd1 vccd1 vccd1 net486
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 team_10_WB.instance_to_wrap.host_row1\[76\] vssd1 vssd1 vccd1 vccd1 net519
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_10_WB.instance_to_wrap.dispFSM.guesses\[5\] vssd1 vssd1 vccd1 vccd1 net530
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold52 team_10_WB.instance_to_wrap.host_row1\[55\] vssd1 vssd1 vccd1 vccd1 net508
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold96 team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs vssd1 vssd1 vccd1 vccd1 net552
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[7\] vssd1 vssd1 vccd1 vccd1
+ net541 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2267__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4014__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3927__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4164__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3240_ net468 _1642_ _1612_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__a21oi_1
X_3171_ _1550_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2122_ net218 net217 team_10_WB.instance_to_wrap.gamelogic.state\[2\] team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__or4b_2
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3455__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2258__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2258__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2053_ team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] net110 net138 net671 vssd1
+ vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2955_ _0798_ _1478_ _0873_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[7\] sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1906_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _0829_ sky130_fd_sc_hd__inv_2
X_2886_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] net1 _1467_ vssd1 vssd1 vccd1
+ vccd1 _1468_ sky130_fd_sc_hd__mux2_1
X_4625_ team_10_WB.instance_to_wrap.lcdPlayer.lcd_en vssd1 vssd1 vccd1 vccd1 net77
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3048__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4556_ net367 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__2194__B1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3507_ net238 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__inv_2
X_4487_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[44\]
+ _0470_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_3438_ _1719_ _1801_ _1810_ net179 vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__a22o_1
X_3369_ team_10_WB.instance_to_wrap.host_row1\[50\] _1699_ net167 team_10_WB.instance_to_wrap.host_row2\[74\]
+ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2249__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3446__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4037__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4187__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3382__C1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1999__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2740_ team_10_WB.instance_to_wrap.clock_div.count\[13\] team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ team_10_WB.instance_to_wrap.clock_div.count\[15\] _1362_ vssd1 vssd1 vccd1 vccd1
+ _1365_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2671_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] _1324_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__o21ai_1
X_4410_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[7\]
+ _0393_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4341_ clknet_leaf_16_wb_clk_i _0731_ _0330_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[64\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4272_ clknet_leaf_0_wb_clk_i _0662_ _0261_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_185_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3223_ net172 _1631_ _1632_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__nor3_1
XFILLER_0_185_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3154_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\] _0899_ _1582_ vssd1
+ vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__or3b_1
X_4569__444 vssd1 vssd1 vccd1 vccd1 net444 _4569__444/LO sky130_fd_sc_hd__conb_1
XANTENNA__3428__B1 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2105_ team_10_WB.instance_to_wrap.dispFSM.guesses\[15\] net144 net108 net482 vssd1
+ vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a22o_1
X_3085_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__mux2_1
X_2036_ team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] net110 net135 team_10_WB.instance_to_wrap.dispFSM.msg\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3987_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[24\]
+ _0055_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2938_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\] net152 net124 net652 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[43\] sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_28_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4541__352 vssd1 vssd1 vccd1 vccd1 _4541__352/HI net352 sky130_fd_sc_hd__conb_1
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2190__B team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2869_ net719 net158 _1302_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.next_state
+ sky130_fd_sc_hd__a21o_1
X_4608_ net382 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4539_ net350 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_159_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3355__C1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3370__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4202__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3940__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4352__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3910_ net289 vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__inv_2
X_4525__336 vssd1 vssd1 vccd1 vccd1 _4525__336/HI net336 sky130_fd_sc_hd__conb_1
X_3841_ net271 vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3772_ net293 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2291__A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2723_ net692 _1354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[8\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2654_ _1228_ _1309_ _1315_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
X_2585_ _1265_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__and2_1
X_4324_ clknet_leaf_21_wb_clk_i net569 _0313_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3361__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout117 _0875_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
Xfanout128 _1188_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
X_4255_ clknet_leaf_6_wb_clk_i _0649_ _0244_ vssd1 vssd1 vccd1 vccd1 team_10_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
Xfanout139 net142 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_3206_ _1621_ _1611_ _1620_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__and3b_1
X_4186_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[48\]
+ _0175_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[48\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4612__386 vssd1 vssd1 vccd1 vccd1 _4612__386/HI net386 sky130_fd_sc_hd__conb_1
XANTENNA__3061__S net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3137_ _1275_ _1550_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__or2_1
X_3068_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] _1528_ net208 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[70\] sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2019_ _0890_ net227 net221 vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout158_X net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2927__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2388__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4225__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\] vssd1 vssd1 vccd1
+ vccd1 net616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3352__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold171 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\] vssd1 vssd1 vccd1 vccd1
+ net627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] vssd1 vssd1 vccd1 vccd1
+ net649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\] vssd1 vssd1 vccd1
+ vccd1 net638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4375__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4364__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3343__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2370_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__a21o_1
X_4040_ clknet_leaf_21_wb_clk_i _0525_ _0081_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4274__Q team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4248__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3824_ net252 vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3755_ net261 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2706_ net607 net536 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3686_ net251 vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_154_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout118_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2637_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _1085_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ _1303_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a221o_1
XANTENNA__4398__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2568_ _0974_ _1253_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__nor2_1
X_4307_ clknet_leaf_15_wb_clk_i _0697_ _0296_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[30\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_113_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2499_ net220 _1218_ _1217_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__mux2_1
X_4238_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[2\]
+ _0227_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3098__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4169_ clknet_leaf_2_wb_clk_i _0638_ _0158_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3325__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3490__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1870_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] vssd1 vssd1 vccd1 vccd1
+ _0795_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3665__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3540_ net245 vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3471_ team_10_WB.instance_to_wrap.dispFSM.guesses\[63\] net173 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[15\]
+ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2422_ net159 net157 vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__nand2_1
X_2353_ _1099_ _1124_ _1125_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__or3_1
XANTENNA__4269__Q team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4023_ clknet_leaf_0_wb_clk_i net485 _0070_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2284_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _1065_ vssd1 vssd1 vccd1
+ vccd1 _1066_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4683__435 vssd1 vssd1 vccd1 vccd1 _4683__435/HI net435 sky130_fd_sc_hd__conb_1
XFILLER_0_126_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3807_ net278 vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1999_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] net147 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1 vccd1 vccd1 _0750_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_115_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3738_ net284 vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__inv_2
X_3669_ net267 vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4413__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2046__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3467__D1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4093__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3482__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\] _0834_ net161 vssd1 vssd1 vccd1
+ vccd1 _1486_ sky130_fd_sc_hd__a41o_1
XFILLER_0_173_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1922_ net299 net5 vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__and2b_1
X_4641_ net409 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_71_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4572_ net447 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3523_ net232 vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__inv_2
X_3454_ team_10_WB.instance_to_wrap.host_row1\[70\] _1703_ net179 team_10_WB.instance_to_wrap.host_row2\[70\]
+ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2405_ team_10_WB.instance_to_wrap.clock_div.count\[14\] team_10_WB.instance_to_wrap.clock_div.count\[17\]
+ team_10_WB.instance_to_wrap.clock_div.count\[16\] team_10_WB.instance_to_wrap.clock_div.count\[15\]
+ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__or4bb_1
X_3385_ team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] net171 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__a22o_1
XANTENNA__4436__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2336_ _1103_ _1104_ _1105_ _1106_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__and4_1
XANTENNA__2458__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2267_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] _0801_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout185_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4006_ clknet_leaf_27_wb_clk_i _0494_ net241 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2276__A2 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2198_ _0976_ _0977_ _0980_ _0985_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2433__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold31 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[1\] vssd1 vssd1
+ vccd1 vccd1 net476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_10_WB.instance_to_wrap.host_row1\[47\] vssd1 vssd1 vccd1 vccd1 net498
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_10_WB.instance_to_wrap.message_reg.msg\[0\] vssd1 vssd1 vccd1 vccd1 net520
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _0591_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 _0672_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] vssd1 vssd1 vccd1
+ vccd1 net553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[7\] vssd1 vssd1 vccd1
+ vccd1 net542 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4372__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3953__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3419__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4309__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4459__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3170_ _0903_ _1277_ net195 vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__and3b_1
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2121_ team_10_WB.instance_to_wrap.gamelogic.state\[2\] _0923_ team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__and3b_1
X_2052_ team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] net110 net138 net701 vssd1
+ vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2954_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\] net163 _1478_ team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[6\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1905_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _0828_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2885_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] vssd1 vssd1 vccd1 vccd1
+ _1467_ sky130_fd_sc_hd__and3b_1
XFILLER_0_154_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4624_ net393 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4555_ net366 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_114_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3391__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3506_ net232 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__inv_2
X_4486_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[43\]
+ _0469_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3064__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3437_ _1799_ _1803_ _1808_ _1811_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__or4_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3368_ net479 net177 _1746_ net229 vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__o211a_1
XANTENNA__2188__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2319_ _0867_ _1090_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__or2_1
X_3299_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout188_X net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3976__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2957__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4367__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4131__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2670_ _1324_ _1325_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4281__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3373__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1923__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4340_ clknet_leaf_22_wb_clk_i _0730_ _0329_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_4271_ clknet_leaf_0_wb_clk_i _0661_ _0260_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3222_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ _1628_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__and3_1
X_3153_ net220 net221 net226 vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__o21a_1
XANTENNA__3999__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2104_ team_10_WB.instance_to_wrap.dispFSM.guesses\[8\] net115 net140 net712 vssd1
+ vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__o22a_1
X_3084_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] _1536_ net208 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[78\] sky130_fd_sc_hd__mux2_1
X_2035_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] net144 net107 net614 vssd1 vssd1
+ vccd1 vccd1 _0744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout148_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3986_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[23\]
+ _0054_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2937_ net215 net151 net120 net685 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[42\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3059__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2868_ net492 _1455_ net176 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[10\]
+ sky130_fd_sc_hd__o21a_1
X_4607_ net381 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__4679__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2799_ _1407_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__inv_2
X_4538_ net349 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4469_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[26\]
+ _0452_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4154__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3310__D_N net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3840_ net267 vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3771_ net261 vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2722_ _1180_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[7\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_124_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2653_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] _0827_ _1225_ _1233_
+ _1313_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__o221a_1
X_2584_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__inv_2
X_4323_ clknet_leaf_15_wb_clk_i _0713_ _0312_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[46\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_2
Xfanout129 _1184_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
Xfanout107 net108 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_2
X_4254_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[10\]
+ _0243_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3205_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] _1392_ vssd1 vssd1 vccd1 vccd1
+ _1621_ sky130_fd_sc_hd__and4_1
XANTENNA__4177__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4185_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[47\]
+ _0174_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[47\] sky130_fd_sc_hd__dfrtp_1
X_3136_ _0903_ _1566_ _1280_ _1277_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__o211a_1
X_3067_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2018_ _0892_ net231 net2 vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__or3b_1
XFILLER_0_54_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3969_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[6\]
+ _0037_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold150 team_10_WB.instance_to_wrap.host_row1\[70\] vssd1 vssd1 vccd1 vccd1 net606
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold161 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\] vssd1 vssd1 vccd1 vccd1
+ net617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] vssd1 vssd1 vccd1 vccd1
+ net639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] vssd1 vssd1 vccd1 vccd1
+ net650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] vssd1 vssd1 vccd1 vccd1
+ net628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4548__359 vssd1 vssd1 vccd1 vccd1 _4548__359/HI net359 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_177_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4380__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3427__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2000__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_184_Right_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3823_ net287 vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__inv_2
XANTENNA__3016__C1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_3754_ net283 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2705_ net536 _1171_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[0\]
+ sky130_fd_sc_hd__nor2_1
X_3685_ net250 vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_154_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2636_ net166 _1301_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_65_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4653__421 vssd1 vssd1 vccd1 vccd1 _4653__421/HI net421 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2567_ _1047_ _1252_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1
+ vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2498_ _0812_ _0888_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__nor2_1
X_4306_ clknet_leaf_21_wb_clk_i _0696_ _0295_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_4237_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[1\]
+ _0226_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4168_ clknet_leaf_29_wb_clk_i _0637_ _0157_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_65_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4099_ clknet_leaf_12_wb_clk_i _0570_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout170_X net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3119_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1278_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_66_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3022__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_83_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4342__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4492__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4637__405 vssd1 vssd1 vccd1 vccd1 _4637__405/HI net405 sky130_fd_sc_hd__conb_1
XFILLER_0_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3470_ team_10_WB.instance_to_wrap.dispFSM.guesses\[23\] net174 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3681__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2421_ net163 net152 vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__nor2_2
X_2352_ _1117_ _1122_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__and3_1
XANTENNA__2524__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2283_ team_10_WB.instance_to_wrap.gamelogic.rights\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4022_ clknet_leaf_0_wb_clk_i net599 _0069_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4215__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3806_ net283 vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout130_A _1183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4365__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3737_ net283 vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__inv_2
X_1998_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] net147 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1 vccd1 _0751_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3668_ net291 vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__inv_2
XANTENNA__4687__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3599_ net282 vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2619_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_183_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2451__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_X clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout290 net298 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_77_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3482__A2 _1854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload6_A clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4388__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2970_ _0835_ net161 vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__nor2_1
XANTENNA__2442__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1921_ net299 net4 vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__and2b_1
XFILLER_0_173_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4640_ net408 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__2993__B2 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4571_ net446 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
X_3522_ net232 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_139_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3453_ team_10_WB.instance_to_wrap.host_row2\[86\] _1686_ _1695_ net303 vssd1 vssd1
+ vccd1 vccd1 _1827_ sky130_fd_sc_hd__a31o_1
X_2404_ _1165_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__or2_1
X_3384_ net465 net177 _1761_ net229 vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_110_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2335_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\] _1089_ vssd1 vssd1
+ vccd1 vccd1 _1111_ sky130_fd_sc_hd__xnor2_1
X_2266_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] net216 vssd1 vssd1 vccd1
+ vccd1 _1048_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_162_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4005_ clknet_leaf_27_wb_clk_i _0493_ net244 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2197_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] net211 vssd1 vssd1 vccd1
+ vccd1 _0986_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout178_A _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3473__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_148_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2433__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_157_Left_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3161__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold32 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] vssd1 vssd1 vccd1 vccd1
+ net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net67 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_10_WB.instance_to_wrap.message_reg.state\[1\] vssd1 vssd1 vccd1 vccd1
+ net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_10_WB.instance_to_wrap.host_row1\[40\] vssd1 vssd1 vccd1 vccd1 net510
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_10_WB.instance_to_wrap.host_row1\[41\] vssd1 vssd1 vccd1 vccd1 net499
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 team_10_WB.instance_to_wrap.host_row1\[65\] vssd1 vssd1 vccd1 vccd1 net554
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold87 team_10_WB.instance_to_wrap.host_row1\[50\] vssd1 vssd1 vccd1 vccd1 net543
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\] vssd1 vssd1 vccd1
+ vccd1 net532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_166_Left_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2975__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3435__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4060__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2120_ net218 net217 vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__nor2_1
X_2051_ net741 net143 net108 net564 vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a22o_1
XANTENNA__3455__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2953_ _0800_ _1478_ _1474_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[5\]
+ sky130_fd_sc_hd__o21ai_1
X_1904_ net290 vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2884_ _1222_ _1466_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[4\]
+ sky130_fd_sc_hd__and2_1
X_4623_ team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs vssd1 vssd1 vccd1 vccd1 net76
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4554_ net365 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_114_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4403__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3505_ net238 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4485_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[42\]
+ _0468_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkload32_A clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3436_ _1715_ _1720_ net231 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1
+ vccd1 vccd1 _1811_ sky130_fd_sc_hd__o211a_1
X_3367_ net179 _1744_ _1745_ _1743_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2318_ team_10_WB.instance_to_wrap.host_col\[3\] _0868_ _1092_ net228 _0856_ vssd1
+ vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o311ai_1
X_3298_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__nor2_1
XANTENNA__3080__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2249_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] _0799_ net213 _0794_ _1030_
+ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__a221o_1
XANTENNA__3446__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3382__B2 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4592__455 vssd1 vssd1 vccd1 vccd1 net455 _4592__455/LO sky130_fd_sc_hd__conb_1
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XANTENNA_input23_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1999__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2948__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3070__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4426__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1923__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4270_ clknet_leaf_2_wb_clk_i _0660_ _0259_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3221_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ net633 vssd1
+ vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3152_ team_10_WB.instance_to_wrap.dispFSM.msg\[2\] _1290_ _1550_ _1283_ vssd1 vssd1
+ vccd1 vccd1 _1581_ sky130_fd_sc_hd__o31a_1
X_2103_ team_10_WB.instance_to_wrap.dispFSM.guesses\[9\] net109 net135 net634 vssd1
+ vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1921__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3083_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__mux2_1
XANTENNA__3428__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2034_ team_10_WB.instance_to_wrap.dispFSM.guesses\[78\] net112 net141 team_10_WB.instance_to_wrap.dispFSM.msg\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2939__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3985_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[22\]
+ _0053_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2936_ net216 net154 net122 net698 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[41\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2867_ _1455_ _1456_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[9\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_157_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4606_ net380 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
X_2798_ _0815_ net178 _1406_ net293 vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__a211o_2
X_4537_ net348 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XANTENNA__3075__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4468_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[25\]
+ _0451_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\]
+ sky130_fd_sc_hd__dfstp_1
X_3419_ team_10_WB.instance_to_wrap.host_row2\[68\] team_10_WB.instance_to_wrap.dispFSM.guesses\[44\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__mux2_1
XANTENNA__3116__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4399_ clknet_leaf_5_wb_clk_i _0784_ _0382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3104__A team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4449__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3052__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3770_ net284 vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__inv_2
X_2721_ team_10_WB.instance_to_wrap.clock_div.count\[7\] _1351_ vssd1 vssd1 vccd1
+ vccd1 _1354_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2652_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2583_ _1256_ _1258_ _1266_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__or4_1
X_4322_ clknet_leaf_21_wb_clk_i _0712_ _0311_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout119 _0875_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_4
X_4253_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[9\]
+ _0242_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout108 _0915_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
X_3204_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\] _1619_ vssd1 vssd1 vccd1
+ vccd1 _1620_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1932__A team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4184_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[46\]
+ _0173_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[46\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3135_ _1561_ _1565_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__xnor2_1
X_3066_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _1527_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[69\] sky130_fd_sc_hd__mux2_1
X_2017_ net2 net300 _0893_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout160_A _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2482__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3968_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[5\]
+ _0036_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3034__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2919_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\] net155 net123 net659
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[24\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_118_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3899_ net255 vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold162 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 team_10_WB.instance_to_wrap.clock_div.count\[1\] vssd1 vssd1 vccd1 vccd1
+ net607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 net596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 team_10_WB.instance_to_wrap.dispFSM.guesses\[75\] vssd1 vssd1 vccd1 vccd1
+ net640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] vssd1 vssd1 vccd1 vccd1
+ net651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4121__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3025__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3989__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3009__A team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2000__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2000__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4531__342 vssd1 vssd1 vccd1 vccd1 _4531__342/HI net342 sky130_fd_sc_hd__conb_1
XFILLER_0_188_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_111_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3822_ net273 vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3753_ net283 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2704_ team_10_WB.instance_to_wrap.host_col\[3\] team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\]
+ net300 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__mux2_1
X_3684_ net245 vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_120_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2635_ _0841_ _1086_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__nor2_2
XANTENNA__4144__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4305_ clknet_leaf_18_wb_clk_i _0695_ _0294_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_2566_ net217 _0948_ _0919_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2497_ net219 _0891_ _1217_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4294__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4236_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[0\]
+ _0225_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4167_ clknet_leaf_29_wb_clk_i _0636_ _0156_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3098__A3 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3118_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] _1278_ vssd1 vssd1 vccd1 vccd1
+ _1549_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4098_ clknet_leaf_12_wb_clk_i _0569_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_66_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3049_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4515__326 vssd1 vssd1 vccd1 vccd1 _4515__326/HI net326 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_6_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4017__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3011__B net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4167__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4602__376 vssd1 vssd1 vccd1 vccd1 _4602__376/HI net376 sky130_fd_sc_hd__conb_1
XANTENNA__1980__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2420_ net204 _0942_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2351_ _1094_ _1097_ net224 _0869_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__o2bb2a_1
X_2282_ _0990_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4021_ clknet_leaf_0_wb_clk_i net556 _0068_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3348__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1997_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] net147 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1 vccd1 vccd1 _0752_
+ sky130_fd_sc_hd__o22a_1
X_3805_ net262 vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3736_ net262 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1971__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3667_ net286 vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3598_ net277 vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2618_ _1294_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] _1074_ vssd1 vssd1
+ vccd1 vccd1 _0006_ sky130_fd_sc_hd__mux2_1
XANTENNA__3083__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2549_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\]
+ _1240_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\] vssd1 vssd1
+ vccd1 vccd1 _1241_ sky130_fd_sc_hd__o31a_2
X_4219_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[81\]
+ _0208_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[81\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3476__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4386__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout291 net294 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_4
Xfanout280 net285 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1920_ net299 net2 vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__and2b_1
XANTENNA__2993__A2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4570_ net445 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_114_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3521_ net232 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2800__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3452_ team_10_WB.instance_to_wrap.host_row1\[54\] _1699_ net181 team_10_WB.instance_to_wrap.host_row2\[62\]
+ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__a22o_1
X_3383_ net302 _1758_ _1759_ net169 _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__a221o_1
X_2403_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ team_10_WB.instance_to_wrap.clock_div.count\[25\] team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__or4_1
XANTENNA__1924__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2334_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\] _0868_ vssd1 vssd1
+ vccd1 vccd1 _1110_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_110_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3458__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2265_ _1035_ _1040_ _1046_ _0949_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__a31o_1
XANTENNA__1940__A team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2196_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _0801_ _0978_ _0979_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__a221o_1
X_4004_ clknet_leaf_27_wb_clk_i _0492_ net241 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2130__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4332__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1939__X _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout240_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4482__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3078__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3719_ net251 vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
Xhold22 team_10_WB.instance_to_wrap.host_row1\[62\] vssd1 vssd1 vccd1 vccd1 net478
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 team_10_WB.instance_to_wrap.host_row1\[61\] vssd1 vssd1 vccd1 vccd1 net467
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 team_10_WB.instance_to_wrap.host_row1\[73\] vssd1 vssd1 vccd1 vccd1 net500
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 team_10_WB.instance_to_wrap.host_row1\[44\] vssd1 vssd1 vccd1 vccd1 net511
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3449__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 team_10_WB.instance_to_wrap.message_reg.msg\[1\] vssd1 vssd1 vccd1 vccd1 net489
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_10_WB.instance_to_wrap.clock_div.count\[6\] vssd1 vssd1 vccd1 vccd1 net533
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] vssd1 vssd1 vccd1
+ vccd1 net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] vssd1 vssd1 vccd1
+ vccd1 net522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] vssd1 vssd1 vccd1 vccd1 net555
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4205__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4355__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2050_ team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] net115 net140 net708 vssd1
+ vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_179_Right_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2952_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] net163 _1478_ net213 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[4\] sky130_fd_sc_hd__o22a_1
XANTENNA__2415__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4608__382 vssd1 vssd1 vccd1 vccd1 _4608__382/HI net382 sky130_fd_sc_hd__conb_1
XFILLER_0_32_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1903_ team_10_WB.instance_to_wrap.uart_receiver.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _0827_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2883_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] _1465_ vssd1 vssd1 vccd1
+ vccd1 _1466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4622_ team_10_WB.instance_to_wrap.uart_transmitter.tx_serial vssd1 vssd1 vccd1 vccd1
+ net75 sky130_fd_sc_hd__clkbuf_1
X_4553_ net364 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4484_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[41\]
+ _0467_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3391__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3504_ net238 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2530__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3435_ team_10_WB.instance_to_wrap.host_row2\[69\] team_10_WB.instance_to_wrap.dispFSM.guesses\[45\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3366_ net209 _0817_ _1690_ _1403_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3297_ net497 _1677_ _1678_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout190_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2317_ net228 _0848_ net196 team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1
+ vccd1 vccd1 _1093_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout288_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2248_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] _0801_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2179_ team_10_WB.instance_to_wrap.correct\[0\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XANTENNA__4378__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3300__A team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3373__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2203__X _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3220_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ _1630_ vssd1
+ vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3151_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] _1551_ _1579_ _1580_ vssd1 vssd1
+ vccd1 vccd1 _0497_ sky130_fd_sc_hd__o22a_1
X_2102_ team_10_WB.instance_to_wrap.dispFSM.guesses\[10\] net111 net136 net626 vssd1
+ vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3082_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _1535_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[77\] sky130_fd_sc_hd__mux2_1
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] net145 net107 net585 vssd1 vssd1
+ vccd1 vccd1 _0746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_185_Left_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3984_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[21\]
+ _0052_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2935_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] net155 net123 net730 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[40\] sky130_fd_sc_hd__o22a_1
XFILLER_0_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2866_ net734 _1454_ net176 vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4605_ net379 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_2797_ team_10_WB.instance_to_wrap.lcdPlayer.currentState\[3\] net178 vssd1 vssd1
+ vccd1 vccd1 _1406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4536_ net347 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout203_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4467_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[24\]
+ _0450_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_4398_ clknet_leaf_6_wb_clk_i _0783_ _0381_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[35\]
+ sky130_fd_sc_hd__dfstp_1
X_3418_ _1790_ _1793_ net302 vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__o21a_1
XANTENNA_input8_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ _1680_ _1718_ net179 _1728_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_168_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2943__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4050__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3355__A2 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4394__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2094__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2720_ team_10_WB.instance_to_wrap.clock_div.count\[7\] _1351_ vssd1 vssd1 vccd1
+ vccd1 _1353_ sky130_fd_sc_hd__or2_1
X_2651_ _1310_ _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2582_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] _1259_ _0901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__a2bb2o_1
X_4321_ clknet_leaf_19_wb_clk_i _0711_ _0310_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[44\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout109 net116 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
X_4252_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[8\]
+ _0241_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3203_ _1619_ _1611_ _1618_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__and3b_1
XFILLER_0_129_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4183_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[45\]
+ _0172_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[45\] sky130_fd_sc_hd__dfrtp_1
X_3134_ _1563_ _1564_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] _0906_
+ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_145_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3065_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__mux2_1
X_2016_ net4 _0887_ _0892_ net227 vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__or4b_2
XFILLER_0_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3967_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[4\]
+ _0035_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2918_ net620 net156 net125 net643 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[23\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3898_ net273 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2849_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\] _1442_ vssd1 vssd1
+ vccd1 vccd1 _1445_ sky130_fd_sc_hd__or2_1
X_4519_ net330 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold152 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\] vssd1 vssd1 vccd1
+ vccd1 net608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\] vssd1 vssd1 vccd1
+ vccd1 net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 team_10_WB.instance_to_wrap.dispFSM.guesses\[71\] vssd1 vssd1 vccd1 vccd1
+ net597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\] vssd1 vssd1 vccd1
+ vccd1 net630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 team_10_WB.instance_to_wrap.clock_div.count\[28\] vssd1 vssd1 vccd1 vccd1
+ net619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\] vssd1 vssd1 vccd1
+ vccd1 net641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] vssd1 vssd1 vccd1
+ vccd1 net652 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4416__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4628__396 vssd1 vssd1 vccd1 vccd1 _4628__396/HI net396 sky130_fd_sc_hd__conb_1
XFILLER_0_138_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2000__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4096__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3821_ net247 vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3752_ net278 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3683_ net283 vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2703_ team_10_WB.instance_to_wrap.host_col\[2\] net220 net300 vssd1 vssd1 vccd1
+ vccd1 net80 sky130_fd_sc_hd__mux2_1
XFILLER_0_112_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2634_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ _1083_ _1075_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__o31a_1
X_2565_ _0974_ _1251_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nor2_1
X_4304_ clknet_leaf_16_wb_clk_i _0694_ _0293_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[27\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_113_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4439__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2496_ net226 _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__nor2_2
X_4235_ clknet_leaf_22_wb_clk_i _0648_ _0224_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_156_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4166_ clknet_leaf_30_wb_clk_i _0635_ _0155_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3117_ net638 net5 _1548_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4097_ clknet_leaf_12_wb_clk_i _0568_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout270_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3048_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _1518_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[60\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4554__365 vssd1 vssd1 vccd1 vccd1 _4554__365/HI net365 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_6_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1980__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1980__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2350_ _1124_ _1125_ _1099_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__o21ai_1
X_2281_ _1012_ _1061_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__or3_2
X_4020_ clknet_leaf_0_wb_clk_i net516 _0067_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2460__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4111__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3804_ net284 vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2533__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1996_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _0874_ _0884_ net158 vssd1
+ vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__o211a_1
X_4497__308 vssd1 vssd1 vccd1 vccd1 _4497__308/HI net308 sky130_fd_sc_hd__conb_1
XFILLER_0_144_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3735_ net279 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1971__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1971__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3666_ net259 vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__inv_2
X_4538__349 vssd1 vssd1 vccd1 vccd1 _4538__349/HI net349 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_171_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3597_ net281 vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2617_ _0830_ _1116_ _1119_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__nor3_1
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2548_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4218_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[80\]
+ _0207_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[80\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2479_ team_10_WB.instance_to_wrap.host_row1\[52\] net130 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__a22o_1
XANTENNA__3979__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4149_ clknet_leaf_17_wb_clk_i _0620_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload0 clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2911__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout292 net294 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_4
XANTENNA__3467__A1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 net285 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_4
Xfanout270 net275 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_77_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4134__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4643__411 vssd1 vssd1 vccd1 vccd1 _4643__411/HI net411 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_103_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2442__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4284__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3520_ net233 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3451_ net592 net177 _1825_ net229 vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__o211a_1
X_3382_ net209 _1690_ _1752_ net231 _1403_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__a221o_1
X_2402_ team_10_WB.instance_to_wrap.clock_div.count\[27\] team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ team_10_WB.instance_to_wrap.clock_div.count\[29\] team_10_WB.instance_to_wrap.clock_div.count\[28\]
+ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__or4_1
X_2333_ _0810_ _0843_ net196 vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__nand3_1
XFILLER_0_137_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2264_ _1038_ _1039_ _1041_ _1043_ _1045_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__a2111oi_1
X_2195_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _0802_ _0981_ _0983_ vssd1
+ vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__o211a_1
X_4003_ clknet_leaf_27_wb_clk_i _0491_ net241 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1979_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net147 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout119_X net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3718_ net250 vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__inv_2
X_3649_ net287 vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4007__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\] vssd1 vssd1 vccd1 vccd1
+ net468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 net65 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2011__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold56 team_10_WB.instance_to_wrap.host_row1\[71\] vssd1 vssd1 vccd1 vccd1 net512
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 team_10_WB.instance_to_wrap.host_row1\[45\] vssd1 vssd1 vccd1 vccd1 net490
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 team_10_WB.instance_to_wrap.host_row1\[79\] vssd1 vssd1 vccd1 vccd1 net501
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 team_10_WB.instance_to_wrap.host_row1\[43\] vssd1 vssd1 vccd1 vccd1 net545
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4157__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] vssd1 vssd1 vccd1 vccd1 net523
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_191_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3385__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2575__C net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2951_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] net163 _1478_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[3\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__1919__C team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1902_ net204 vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4621_ net392 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2882_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] net223 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__or3b_1
XFILLER_0_154_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3376__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552_ net363 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4483_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[40\]
+ _0466_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\]
+ sky130_fd_sc_hd__dfstp_1
X_3503_ net238 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__inv_2
X_3434_ team_10_WB.instance_to_wrap.host_row2\[85\] team_10_WB.instance_to_wrap.dispFSM.guesses\[61\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3365_ team_10_WB.instance_to_wrap.host_row2\[65\] team_10_WB.instance_to_wrap.dispFSM.guesses\[41\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload18_A clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3296_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ _1674_ net296 vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2316_ net224 net225 _0850_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__and3b_1
X_2247_ _0793_ net212 _0802_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] _1028_
+ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout183_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2178_ _0968_ team_10_WB.instance_to_wrap.correct\[1\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2006__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3118__A team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XANTENNA__4010__Q team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_168_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3300__B _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3358__B1 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4322__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3150_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] _1278_ _1568_ vssd1 vssd1 vccd1
+ vccd1 _1580_ sky130_fd_sc_hd__a21o_1
X_2101_ team_10_WB.instance_to_wrap.dispFSM.guesses\[11\] net113 net139 net715 vssd1
+ vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4472__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3081_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2032_ _0885_ _0903_ net137 vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3983_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[20\]
+ _0051_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2934_ net631 net156 net125 net641 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[39\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2865_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] _1454_ vssd1 vssd1
+ vccd1 vccd1 _1455_ sky130_fd_sc_hd__and2_1
X_4604_ net378 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__3349__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4535_ net346 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2796_ _1405_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4466_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[23\]
+ _0449_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3417_ team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] _1715_ _1791_ _1792_ vssd1
+ vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__a211o_1
X_4397_ clknet_leaf_5_wb_clk_i _0782_ _0380_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[34\]
+ sky130_fd_sc_hd__dfstp_1
X_3348_ team_10_WB.instance_to_wrap.host_row2\[64\] team_10_WB.instance_to_wrap.dispFSM.guesses\[40\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3279_ net593 _1664_ net230 vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2017__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4345__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_X clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_186_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2251__B1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2650_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ _1224_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__or4_1
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2581_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\] _0904_ _0906_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__a22o_1
X_4320_ clknet_leaf_17_wb_clk_i _0710_ _0309_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[43\]
+ sky130_fd_sc_hd__dfstp_1
X_4251_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[7\]
+ _0240_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3202_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\]
+ _1392_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1932__C team_10_WB.instance_to_wrap.host_col\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4182_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[44\]
+ _0171_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[44\] sky130_fd_sc_hd__dfrtp_1
X_3133_ net219 _0905_ _1562_ _0907_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_145_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4218__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3064_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] _1526_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\] sky130_fd_sc_hd__mux2_1
X_2015_ _0887_ _0892_ net227 vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__or3b_1
XANTENNA__2536__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2490__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[3\]
+ _0034_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout146_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4368__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2917_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\] net153 net121 net646
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[22\]
+ sky130_fd_sc_hd__o22a_1
X_3897_ net287 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2848_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\] _1442_ vssd1 vssd1
+ vccd1 vccd1 _1444_ sky130_fd_sc_hd__and2_1
X_2779_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__nand2_1
X_4518_ net329 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xhold153 team_10_WB.instance_to_wrap.host_row1\[54\] vssd1 vssd1 vccd1 vccd1 net609
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 team_10_WB.instance_to_wrap.dispFSM.guesses\[23\] vssd1 vssd1 vccd1 vccd1
+ net587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] vssd1 vssd1 vccd1 vccd1 net598
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[21\] vssd1 vssd1
+ vccd1 vccd1 net576 sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[6\]
+ _0432_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xhold186 team_10_WB.instance_to_wrap.dispFSM.guesses\[14\] vssd1 vssd1 vccd1 vccd1
+ net642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[47\] vssd1 vssd1 vccd1
+ vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\] vssd1 vssd1 vccd1
+ vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 team_10_WB.instance_to_wrap.dispFSM.guesses\[66\] vssd1 vssd1 vccd1 vccd1
+ net653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3016__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3820_ net270 vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_25_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2224__A0 team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3751_ net278 vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2702_ team_10_WB.instance_to_wrap.host_col\[1\] team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\]
+ net300 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__mux2_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3682_ net255 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__inv_2
XANTENNA__1983__C1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2633_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] _1285_ _1290_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1300_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a221o_1
X_2564_ _1059_ _1250_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1
+ vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__a21oi_1
X_4303_ clknet_leaf_17_wb_clk_i _0693_ _0292_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_120_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2495_ net231 _1177_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_34_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4040__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4234_ clknet_leaf_22_wb_clk_i _0647_ _0223_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4165_ clknet_leaf_26_wb_clk_i _0634_ _0154_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3116_ net596 net4 _1548_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__mux2_1
X_4096_ clknet_leaf_12_wb_clk_i _0567_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3047_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__mux2_1
XANTENNA__4190__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4660__428 vssd1 vssd1 vccd1 vccd1 _4660__428/HI net428 sky130_fd_sc_hd__conb_1
XFILLER_0_81_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_176_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3949_ clknet_leaf_23_wb_clk_i _0012_ net256 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4669__431 vssd1 vssd1 vccd1 vccd1 _4669__431/HI net431 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_183_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4565__440 vssd1 vssd1 vccd1 vccd1 net440 _4565__440/LO sky130_fd_sc_hd__conb_1
XFILLER_0_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4063__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2280_ net218 _0952_ _1023_ _1060_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3323__X _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3803_ net261 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1995_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] net146 vssd1 vssd1
+ vccd1 vccd1 _0884_ sky130_fd_sc_hd__or2_1
X_3734_ net292 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__inv_2
X_3665_ net294 vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4406__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1956__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1971__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2616_ _0015_ _0012_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[2\]
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_171_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3596_ net281 vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout109_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2547_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _1239_ sky130_fd_sc_hd__and3b_1
X_2478_ net505 net129 _1189_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__o22a_1
X_4217_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[79\]
+ _0206_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[79\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3476__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4588__451 vssd1 vssd1 vccd1 vccd1 net451 _4588__451/LO sky130_fd_sc_hd__conb_1
X_4148_ clknet_leaf_17_wb_clk_i _0619_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfxtp_1
X_4079_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[10\]
+ _0099_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2009__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2987__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4521__332 vssd1 vssd1 vccd1 vccd1 _4521__332/HI net332 sky130_fd_sc_hd__conb_1
XANTENNA__2025__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload1 clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1864__A team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3164__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 net285 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_77_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2978__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4429__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3465__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3450_ _1781_ _1820_ _1824_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__or3_1
X_2401_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ _1160_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or4_1
X_3381_ team_10_WB.instance_to_wrap.host_row1\[58\] team_10_WB.instance_to_wrap.dispFSM.msg\[2\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__mux2_1
X_2332_ _0843_ net196 _0810_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3458__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2263_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0800_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ _0790_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__a221o_1
X_4002_ clknet_leaf_25_wb_clk_i _0490_ net239 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2194_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _0801_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ _0795_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__o221a_1
XFILLER_0_189_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2969__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2969__B2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4505__316 vssd1 vssd1 vccd1 vccd1 _4505__316/HI net316 sky130_fd_sc_hd__conb_1
XFILLER_0_157_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1978_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] net149 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3717_ net250 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__inv_2
X_3648_ net259 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3579_ net277 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__inv_2
XANTENNA__3946__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 net64 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 _0581_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\] vssd1 vssd1 vccd1 vccd1
+ net480 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] vssd1 vssd1 vccd1
+ vccd1 net513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] vssd1 vssd1 vccd1
+ vccd1 net535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _0509_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4008__Q team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3082__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_193_Right_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4251__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3073__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2950_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\] net164 _1478_ net215 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[2\] sky130_fd_sc_hd__o22a_1
X_1901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _0825_ sky130_fd_sc_hd__inv_2
X_2881_ net193 _1464_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[3\]
+ sky130_fd_sc_hd__and2_1
X_4620_ net391 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4551_ net362 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3969__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3502_ net238 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__inv_2
X_4482_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[39\]
+ _0465_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3433_ team_10_WB.instance_to_wrap.host_row1\[69\] net302 _1703_ vssd1 vssd1 vccd1
+ vccd1 _1808_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3364_ _1738_ _1742_ _1736_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__o21a_1
X_3295_ net296 _1676_ _1677_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__nor3_1
X_2315_ _0868_ _1090_ net4 vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__or3b_1
X_2246_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _0804_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_164_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2177_ _0936_ _0962_ _0967_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3367__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XANTENNA__4124__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__4274__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3055__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2869__B1 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2100_ team_10_WB.instance_to_wrap.dispFSM.guesses\[12\] net113 net139 net658 vssd1
+ vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__o22a_1
X_3080_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] _1534_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[76\] sky130_fd_sc_hd__mux2_1
XFILLER_0_118_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2031_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _0886_ _0910_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_109_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3046__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3982_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[19\]
+ _0050_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_2933_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] net153 net121 net644
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[38\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_150_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2864_ _1454_ net176 _1453_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4603_ net377 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2795_ net230 _1404_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4621__392 vssd1 vssd1 vccd1 vccd1 _4621__392/HI net392 sky130_fd_sc_hd__conb_1
XANTENNA__4147__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4534_ net345 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_159_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4465_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[22\]
+ _0448_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkload30_A clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1962__A team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4396_ clknet_leaf_9_wb_clk_i _0781_ _0379_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4297__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3416_ team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] net171 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[12\]
+ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3347_ _1682_ _1686_ _1688_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_168_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\]
+ _1663_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2229_ net705 net143 _0807_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_127_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3401__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1872__A team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2251__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2251__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2580_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\] _0906_ _1262_ _1263_
+ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__o2111a_1
X_4250_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[6\]
+ _0239_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3201_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\]
+ _1391_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1
+ _1618_ sky130_fd_sc_hd__a31o_1
X_4181_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\]
+ _0170_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[43\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__1932__D team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3132_ _0890_ _0899_ _1259_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__or3_1
XFILLER_0_179_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3063_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2014_ net2 net3 net4 net5 net300 vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__o41a_1
XFILLER_0_54_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3965_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[2\]
+ _0033_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3896_ net269 vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2916_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\] net156 net125 net575
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[21\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout139_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2847_ _1442_ _1443_ net176 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold110 team_10_WB.instance_to_wrap.dispFSM.guesses\[15\] vssd1 vssd1 vccd1 vccd1
+ net566 sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ net461 _1388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[29\]
+ sky130_fd_sc_hd__xor2_1
X_4517_ net328 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
Xhold132 _0690_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _0507_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 team_10_WB.instance_to_wrap.dispFSM.guesses\[13\] vssd1 vssd1 vccd1 vccd1
+ net577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\] vssd1 vssd1 vccd1 vccd1
+ net610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[31\] vssd1 vssd1
+ vccd1 vccd1 net621 sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ clknet_leaf_28_wb_clk_i net481 _0431_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold198 team_10_WB.instance_to_wrap.dispFSM.guesses\[64\] vssd1 vssd1 vccd1 vccd1
+ net654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\] vssd1 vssd1 vccd1
+ vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4379_ clknet_leaf_6_wb_clk_i _0764_ _0362_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_44_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4312__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2481__A1 team_10_WB.instance_to_wrap.host_row1\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2233__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4462__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3750_ net293 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2701_ team_10_WB.instance_to_wrap.host_col\[0\] net222 net300 vssd1 vssd1 vccd1
+ vccd1 net78 sky130_fd_sc_hd__mux2_1
XFILLER_0_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3681_ net294 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2632_ net195 _1281_ _1298_ _0903_ _1299_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__a221o_1
X_2563_ net218 _0948_ _0919_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__o21ai_1
X_4302_ clknet_leaf_18_wb_clk_i _0692_ _0291_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[25\]
+ sky130_fd_sc_hd__dfstp_1
X_2494_ net510 net132 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] vssd1
+ vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__a22o_1
X_4233_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[2\]
+ _0222_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4164_ clknet_leaf_29_wb_clk_i _0633_ _0153_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4095_ clknet_leaf_12_wb_clk_i _0566_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3115_ net571 net3 _1548_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3046_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _1517_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[59\] sky130_fd_sc_hd__mux2_1
XANTENNA__4335__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2463__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2463__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4485__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_176_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3412__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3948_ clknet_leaf_21_wb_clk_i _0011_ net256 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3879_ net277 vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2789__Y _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4208__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4358__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3802_ net280 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1994_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] net147 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1 vccd1 _0754_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3733_ net245 vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3664_ net255 vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload30 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_6
XFILLER_0_42_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2615_ _1270_ _1282_ _1293_ _1275_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_171_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2131__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3595_ net259 vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2546_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nand2b_1
X_2477_ net609 net132 _1185_ _1212_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__a22o_1
X_4216_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[78\]
+ _0205_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[78\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4147_ clknet_leaf_16_wb_clk_i _0618_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfxtp_1
X_4078_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[9\]
+ _0098_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3029_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\]
+ net192 vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload2 clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinvlp_4
X_4560__371 vssd1 vssd1 vccd1 vccd1 _4560__371/HI net371 sky130_fd_sc_hd__conb_1
XANTENNA__2911__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1880__A team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 net251 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_4
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_4
Xfanout272 net275 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_4
XANTENNA__2124__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout261 net264 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout294 net298 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2978__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4180__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2400_ team_10_WB.instance_to_wrap.clock_div.count\[11\] _1161_ _1162_ team_10_WB.instance_to_wrap.clock_div.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__or4b_1
XFILLER_0_122_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3380_ _1754_ _1755_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__or3_1
X_2331_ _0844_ _0855_ _0809_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__a21o_1
XANTENNA__3481__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2262_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] net215 vssd1 vssd1 vccd1
+ vccd1 _1044_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4001_ clknet_leaf_25_wb_clk_i _0489_ net241 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2193_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] _0804_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2969__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4544__355 vssd1 vssd1 vccd1 vccd1 _4544__355/HI net355 sky130_fd_sc_hd__conb_1
XFILLER_0_172_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1977_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] net150 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1965__A team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3716_ net251 vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3647_ net274 vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3578_ net288 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_132_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2529_ net547 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0512_ sky130_fd_sc_hd__mux2_1
Xhold14 team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] vssd1 vssd1 vccd1 vccd1 net470
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\] vssd1 vssd1 vccd1
+ vccd1 net492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[5\] vssd1 vssd1 vccd1
+ vccd1 net481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_10_WB.instance_to_wrap.message_reg.msg\[7\] vssd1 vssd1 vccd1 vccd1 net503
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_10_WB.instance_to_wrap.host_row1\[49\] vssd1 vssd1 vccd1 vccd1 net525
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[1\] vssd1 vssd1
+ vccd1 vccd1 net514 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_39_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3385__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1875__A team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4528__339 vssd1 vssd1 vccd1 vccd1 _4528__339/HI net339 sky130_fd_sc_hd__conb_1
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1900_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] vssd1 vssd1 vccd1 vccd1
+ _0824_ sky130_fd_sc_hd__inv_2
X_2880_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] net1 _1463_ vssd1 vssd1 vccd1
+ vccd1 _1464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3376__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4550_ net361 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4481_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[38\]
+ _0464_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\]
+ sky130_fd_sc_hd__dfstp_1
X_3501_ net238 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__inv_2
X_3432_ team_10_WB.instance_to_wrap.host_row1\[101\] net302 _1776_ _1806_ vssd1 vssd1
+ vccd1 vccd1 _1807_ sky130_fd_sc_hd__o22a_1
X_3363_ _1739_ _1740_ _1741_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__or3_1
XANTENNA__3064__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3294_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\]
+ _1672_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2314_ net224 net225 _0850_ _0818_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__o211ai_1
X_2245_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _0800_ _0802_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__o221a_1
XANTENNA__4076__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2176_ _0959_ _0960_ _0961_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout169_A _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4679_ net184 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_9_wb_clk_i_X clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4633__401 vssd1 vssd1 vccd1 vccd1 _4633__401/HI net401 sky130_fd_sc_hd__conb_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XANTENNA__4419__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2973__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3358__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2213__B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3309__B team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4099__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ net195 _0903_ net143 vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_178_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2097__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3981_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[18\]
+ _0049_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2932_ net740 net156 net125 net586 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[37\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2863_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\]
+ _1450_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602_ net376 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_154_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2794_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[5\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__mux2_1
X_4533_ net344 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_159_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ clknet_leaf_27_wb_clk_i net576 _0447_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2309__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4395_ clknet_leaf_6_wb_clk_i _0780_ _0378_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[32\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkload23_A clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3415_ team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] net173 net168 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\]
+ _1771_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_90_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3346_ _1722_ _1725_ _1713_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_168_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Left_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3277_ net487 _1661_ _1665_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout286_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2228_ net477 _1011_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _0924_ _0945_ _0951_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__or4_1
XFILLER_0_191_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3401__C net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_179_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_172_Left_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_181_Left_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_186_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4391__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3959__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_190_Left_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2539__A0 team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3200_ net172 _1617_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__nor2_1
X_4180_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[42\]
+ _0169_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[42\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2894__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3131_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] _1259_ vssd1 vssd1
+ vccd1 vccd1 _1562_ sky130_fd_sc_hd__nor2_1
X_3062_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] _1525_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[67\] sky130_fd_sc_hd__mux2_1
X_2013_ net300 net5 vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4114__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3964_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[1\]
+ _0032_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3895_ net296 vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__inv_2
X_2915_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\] net151 net120 net736
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[20\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2846_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2777_ _1387_ _1388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[28\]
+ sky130_fd_sc_hd__nor2_1
Xhold100 _0506_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ net327 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
Xhold133 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\] vssd1 vssd1 vccd1
+ vccd1 net589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _0682_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\] vssd1 vssd1 vccd1
+ vccd1 net600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _0680_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] vssd1 vssd1 vccd1 vccd1
+ net633 sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[4\]
+ _0430_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\]
+ sky130_fd_sc_hd__dfstp_1
Xhold166 team_10_WB.instance_to_wrap.dispFSM.guesses\[44\] vssd1 vssd1 vccd1 vccd1
+ net622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 team_10_WB.instance_to_wrap.dispFSM.guesses\[31\] vssd1 vssd1 vccd1 vccd1
+ net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold188 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\] vssd1 vssd1 vccd1
+ vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 team_10_WB.instance_to_wrap.clock_div.count\[4\] vssd1 vssd1 vccd1 vccd1
+ net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2702__A0 team_10_WB.instance_to_wrap.host_col\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_input6_A gpio_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4378_ clknet_leaf_2_wb_clk_i _0763_ _0361_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3329_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _1682_ _1688_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout191_X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2233__A2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2941__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_188_Right_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4137__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3421__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4287__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2700_ _1342_ _1344_ _1238_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.tx_serial
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3680_ net259 vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2631_ _0911_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2562_ _0919_ _0972_ _1249_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__and3_1
X_4301_ clknet_leaf_15_wb_clk_i _0691_ _0290_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_120_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2493_ net499 net133 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] vssd1
+ vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__a22o_1
X_4232_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[1\]
+ _0221_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4163_ clknet_leaf_26_wb_clk_i _0632_ _0152_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4094_ clknet_leaf_12_wb_clk_i _0565_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3114_ net529 net2 _1548_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3045_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__mux2_1
XANTENNA__2129__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2463__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout151_A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3947_ clknet_leaf_2_wb_clk_i _0479_ _0021_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_176_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1974__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3878_ net269 vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__inv_2
X_2829_ _1411_ _1418_ _1426_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__and3_1
XANTENNA__1974__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2439__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2914__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3801_ net279 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__inv_2
X_1993_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] _0874_ _0883_ net159 vssd1
+ vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_71_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1956__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3732_ net249 vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__inv_2
Xclkload20 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_125_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3663_ net281 vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload31 clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2614_ _0824_ _1287_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3594_ net276 vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4302__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2545_ net227 net457 _1216_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__mux2_1
XANTENNA__2381__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4400__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2476_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] net185 vssd1 vssd1 vccd1
+ vccd1 _1212_ sky130_fd_sc_hd__or2_1
X_4215_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[77\]
+ _0204_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[77\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4146_ clknet_leaf_16_wb_clk_i _0617_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout199_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4452__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_32_wb_clk_i_X clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4077_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[8\]
+ _0097_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3028_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] _1508_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[50\] sky130_fd_sc_hd__mux2_1
XANTENNA__2009__D net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload3 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_190_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout240 net266 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_2
Xfanout273 net275 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_4
Xfanout251 net265 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_4
Xfanout295 net296 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout284 net285 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3388__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4325__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2232__A team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4650__418 vssd1 vssd1 vccd1 vccd1 _4650__418/HI net418 sky130_fd_sc_hd__conb_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] _0819_ _0849_ vssd1
+ vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__or3_1
XANTENNA__4475__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2261_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] _0799_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\]
+ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4000_ clknet_leaf_25_wb_clk_i _0488_ net239 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2192_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _0802_ _0804_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_99_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3379__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1976_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _0874_ _0880_ net158 vssd1
+ vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3715_ net267 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3646_ net291 vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3577_ net277 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2528_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__inv_2
Xhold26 team_10_WB.instance_to_wrap.dispFSM.guesses\[7\] vssd1 vssd1 vccd1 vccd1 net482
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 _0511_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_10_WB.instance_to_wrap.message_reg.msg\[3\] vssd1 vssd1 vccd1 vccd1 net493
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] net197 _1185_
+ _1202_ net130 vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__a221o_1
Xhold48 team_10_WB.instance_to_wrap.host_row1\[72\] vssd1 vssd1 vccd1 vccd1 net504
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] vssd1 vssd1 vccd1 vccd1 net515
+ sky130_fd_sc_hd__dlygate4sd3_1
X_4129_ clknet_leaf_10_wb_clk_i _0600_ _0128_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3992__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4348__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3500_ net238 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__inv_2
X_4480_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[37\]
+ _0463_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_3431_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1805_ _1686_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3362_ team_10_WB.instance_to_wrap.host_row2\[49\] net170 _1708_ team_10_WB.instance_to_wrap.host_row1\[73\]
+ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__a22o_1
X_2313_ net228 _0848_ net196 net224 vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_76_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3293_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\] _1674_ vssd1 vssd1 vccd1
+ vccd1 _1676_ sky130_fd_sc_hd__nor2_1
X_2244_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0798_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__o22a_1
X_4511__322 vssd1 vssd1 vccd1 vccd1 _4511__322/HI net322 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_10_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2175_ _0966_ team_10_WB.instance_to_wrap.correct\[2\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2137__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout231_A _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1959_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] net150 _0875_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\]
+ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4678_ net433 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_160_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3629_ net247 vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__inv_2
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4170__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3460__C1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2263__B1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2318__A1 team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2869__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3980_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[17\]
+ _0048_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2931_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] net151 net120 net667
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[36\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_33_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3451__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4601_ net375 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_127_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2862_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ _1448_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\] vssd1 vssd1 vccd1
+ vccd1 _1453_ sky130_fd_sc_hd__a31o_1
X_2793_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] _1393_ _1395_ _1402_
+ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__or4_4
XFILLER_0_25_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4532_ net343 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
X_4656__424 vssd1 vssd1 vccd1 vccd1 _4656__424/HI net424 sky130_fd_sc_hd__conb_1
X_4463_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[20\]
+ _0446_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3414_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1704_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[68\]
+ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__a221o_1
XANTENNA__2420__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2309__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4043__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4394_ clknet_leaf_2_wb_clk_i _0779_ _0377_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_3345_ _1716_ _1723_ _1724_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__or3_1
XANTENNA_clkload16_A clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3276_ net295 _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2227_ team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] _1009_ _1010_ _0808_
+ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout279_A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4193__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2493__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2158_ net218 net217 _0947_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__a31o_1
XFILLER_0_191_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2089_ team_10_WB.instance_to_wrap.dispFSM.guesses\[31\] net145 net107 net587 vssd1
+ vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_179_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600__456 vssd1 vssd1 vccd1 vccd1 net456 _4600__456/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_99_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2236__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_3__f_wb_clk_i_X clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4066__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3130_ _1286_ _1554_ _1560_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__or3b_1
XANTENNA__2894__B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3061_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2012_ net299 net5 vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__and2_1
XANTENNA__2475__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3963_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[0\]
+ _0031_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2914_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\] net155 net123 net664
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[19\]
+ sky130_fd_sc_hd__o22a_1
X_3894_ net288 vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4409__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2845_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1442_ sky130_fd_sc_hd__and3_1
XANTENNA__1986__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4515_ net326 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2776_ team_10_WB.instance_to_wrap.clock_div.count\[27\] team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ team_10_WB.instance_to_wrap.clock_div.count\[28\] _1384_ vssd1 vssd1 vccd1 vccd1
+ _1388_ sky130_fd_sc_hd__and4_1
Xhold101 team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] vssd1 vssd1 vccd1 vccd1 net557
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2421__Y _1183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold123 team_10_WB.instance_to_wrap.host_row1\[75\] vssd1 vssd1 vccd1 vccd1 net579
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\] vssd1 vssd1 vccd1
+ vccd1 net590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 team_10_WB.instance_to_wrap.dispFSM.guesses\[47\] vssd1 vssd1 vccd1 vccd1
+ net568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold167 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\] vssd1 vssd1 vccd1
+ vccd1 net623 sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[3\]
+ _0429_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2950__B2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold145 team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\] vssd1 vssd1 vccd1 vccd1
+ net601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2150__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold156 _0698_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4377_ clknet_leaf_7_wb_clk_i _0762_ _0360_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\]
+ sky130_fd_sc_hd__dfstp_2
Xhold189 team_10_WB.instance_to_wrap.dispFSM.guesses\[8\] vssd1 vssd1 vccd1 vccd1
+ net645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] vssd1 vssd1 vccd1 vccd1
+ net634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _1697_ _1707_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__nor2_4
XFILLER_0_95_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2702__A1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3259_ net295 _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4089__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2941__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2630_ _0886_ _0909_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__nor2_1
XANTENNA__3337__Y _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2561_ net218 net217 _0947_ _1034_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__a41o_1
X_2492_ net582 net133 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\] vssd1
+ vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__a22o_1
X_4300_ clknet_leaf_18_wb_clk_i net588 _0289_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ clknet_leaf_33_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[0\]
+ _0220_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_49_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4162_ clknet_leaf_27_wb_clk_i _0631_ _0151_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4093_ clknet_leaf_12_wb_clk_i _0564_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3113_ net561 net219 _1548_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3044_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] _1516_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[58\] sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_X clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_179_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2999__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3946_ clknet_leaf_2_wb_clk_i _0478_ _0020_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout144_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3412__A2 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1974__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3877_ net252 vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__inv_2
X_2828_ _1409_ _0513_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4381__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2759_ team_10_WB.instance_to_wrap.clock_div.count\[21\] _1376_ vssd1 vssd1 vccd1
+ vccd1 _1378_ sky130_fd_sc_hd__and2_1
XANTENNA__3949__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4429_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[26\]
+ _0412_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3479__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1894__A team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3167__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4572__447 vssd1 vssd1 vccd1 vccd1 net447 _4572__447/LO sky130_fd_sc_hd__conb_1
XANTENNA__3614__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4254__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3800_ net264 vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3731_ net246 vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__inv_2
X_1992_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] net146 vssd1 vssd1
+ vccd1 vccd1 _0883_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3662_ net273 vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload10 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__bufinv_16
Xclkload21 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_4
XFILLER_0_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2613_ _0016_ _0014_ _0015_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
X_3593_ net260 vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__inv_2
Xclkload32 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2544_ team_10_WB.instance_to_wrap.host_col\[0\] _1237_ _1179_ vssd1 vssd1 vccd1
+ vccd1 _0484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2475_ net508 net130 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__a22o_1
X_4214_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[76\]
+ _0203_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[76\] sky130_fd_sc_hd__dfrtp_1
X_4145_ clknet_leaf_19_wb_clk_i _0616_ _0144_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4076_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[7\]
+ _0096_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3027_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout261_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3929_ net271 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__inv_2
Xclkload4 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_16
XFILLER_0_190_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4127__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 _0018_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
XANTENNA__4277__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout241 net244 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_4
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_4
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_4
Xfanout252 net265 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_4
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout285 net298 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3085__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3328__B _1707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2232__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2899__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2260_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0800_ vssd1 vssd1 vccd1
+ vccd1 _1042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2191_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] team_10_WB.instance_to_wrap.gamelogic.letter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_162_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1975_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] net146 vssd1 vssd1 vccd1
+ vccd1 _0880_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3714_ net250 vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3645_ net270 vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3576_ net274 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2527_ team_10_WB.instance_to_wrap.uart_receiver.state\[0\] team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] vssd1 vssd1 vccd1 vccd1 _1233_
+ sky130_fd_sc_hd__or3b_4
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2458_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] net185 vssd1 vssd1 vccd1
+ vccd1 _1202_ sky130_fd_sc_hd__or2_1
Xhold16 net68 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 _0674_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold38 team_10_WB.instance_to_wrap.message_reg.msg\[2\] vssd1 vssd1 vccd1 vccd1 net494
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_10_WB.instance_to_wrap.host_row1\[53\] vssd1 vssd1 vccd1 vccd1 net505
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _0844_ net570 _1158_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__mux2_1
X_4128_ clknet_leaf_28_wb_clk_i _0599_ _0127_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_4059_ clknet_leaf_14_wb_clk_i _0544_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3067__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input37_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3058__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2805__A0 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3103__S net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2243__A team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4442__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3430_ net209 _0817_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3361_ team_10_WB.instance_to_wrap.host_row1\[49\] _1699_ net169 team_10_WB.instance_to_wrap.host_row1\[57\]
+ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2312_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__inv_2
X_3292_ net488 _1672_ _1675_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3802__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2243_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] _0805_ vssd1 vssd1 vccd1
+ vccd1 _1025_ sky130_fd_sc_hd__or2_1
XANTENNA__3361__X _1740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4550__361 vssd1 vssd1 vccd1 vccd1 _4550__361/HI net361 sky130_fd_sc_hd__conb_1
XFILLER_0_164_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2174_ _0964_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3049__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2424__Y _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1958_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] net148 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[35\]
+ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1889_ net732 vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__inv_2
X_4677_ net183 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3628_ net248 vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__inv_2
X_3559_ net240 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__inv_2
XANTENNA__3288__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4315__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3460__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2263__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4465__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2998__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4493__304 vssd1 vssd1 vccd1 vccd1 _4493__304/HI net304 sky130_fd_sc_hd__conb_1
X_4534__345 vssd1 vssd1 vccd1 vccd1 _4534__345/HI net345 sky130_fd_sc_hd__conb_1
XANTENNA__3279__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4226__Q team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2930_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] net155 net123 net672
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[35\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_33_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4600_ net456 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_0_127_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2861_ net522 _1450_ _1452_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_2792_ _1396_ _1400_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__or3_1
XFILLER_0_127_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4531_ net342 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4462_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[19\]
+ _0445_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3413_ team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] net181 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a22o_1
XANTENNA__3982__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4393_ clknet_leaf_7_wb_clk_i _0778_ _0376_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2420__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3344_ team_10_WB.instance_to_wrap.dispFSM.guesses\[0\] _1717_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[64\]
+ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3275_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] _1661_ vssd1 vssd1 vccd1
+ vccd1 _1664_ sky130_fd_sc_hd__and2_1
X_2226_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _1010_ sky130_fd_sc_hd__or3b_1
XANTENNA__4338__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2157_ net217 _0916_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__nor2_1
X_2088_ team_10_WB.instance_to_wrap.dispFSM.guesses\[24\] net114 net140 net722 vssd1
+ vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_127_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4488__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2245__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2245__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4518__329 vssd1 vssd1 vccd1 vccd1 _4518__329/HI net329 sky130_fd_sc_hd__conb_1
XFILLER_0_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3433__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4605__379 vssd1 vssd1 vccd1 vccd1 _4605__379/HI net379 sky130_fd_sc_hd__conb_1
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3617__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3060_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] _1524_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[66\] sky130_fd_sc_hd__mux2_1
XFILLER_0_173_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_X clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2011_ net299 net4 vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4582__449 vssd1 vssd1 vccd1 vccd1 net449 _4582__449/LO sky130_fd_sc_hd__conb_1
XFILLER_0_161_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3424__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3962_ clknet_leaf_22_wb_clk_i _0482_ _0030_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3893_ net270 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__inv_2
X_2913_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\] net151 net120 net714
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[18\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2844_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] net475 _1441_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4010__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4514_ net325 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__2431__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2775_ team_10_WB.instance_to_wrap.clock_div.count\[27\] _1386_ net619 vssd1 vssd1
+ vccd1 vccd1 _1387_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold135 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\] vssd1 vssd1 vccd1
+ vccd1 net591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _0510_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] vssd1 vssd1 vccd1
+ vccd1 net580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _0714_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold157 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4445_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[2\]
+ _0428_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\]
+ sky130_fd_sc_hd__dfstp_1
Xhold146 team_10_WB.instance_to_wrap.clock_div.count\[24\] vssd1 vssd1 vccd1 vccd1
+ net602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_10_WB.instance_to_wrap.dispFSM.guesses\[63\] vssd1 vssd1 vccd1 vccd1
+ net624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\] vssd1 vssd1 vccd1
+ vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4160__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4376_ clknet_leaf_2_wb_clk_i _0761_ _0359_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_186_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3360__C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3327_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _0817_ vssd1 vssd1 vccd1
+ vccd1 _1707_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout291_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] _1651_ vssd1 vssd1 vccd1
+ vccd1 _1653_ sky130_fd_sc_hd__and2_1
X_3189_ net297 net178 _1610_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2209_ net517 _0996_ _0992_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__o21a_1
XANTENNA__2466__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3415__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1977__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2941__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3351__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3900__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4033__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1968__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4499__310 vssd1 vssd1 vccd1 vccd1 _4499__310/HI net310 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_117_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4183__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ _0973_ _1248_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and2_1
X_2491_ net545 net132 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] vssd1
+ vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4230_ clknet_leaf_1_wb_clk_i _0646_ _0219_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_4161_ clknet_leaf_30_wb_clk_i _0630_ _0150_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4092_ clknet_leaf_8_wb_clk_i _0563_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3112_ net540 net220 _1548_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3043_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3810__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3945_ clknet_leaf_4_wb_clk_i _0477_ _0019_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_147_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1959__B1 _0875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout137_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3876_ net252 vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__inv_2
X_2827_ _1407_ _1418_ _1429_ _1427_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2758_ team_10_WB.instance_to_wrap.clock_div.count\[21\] _1376_ vssd1 vssd1 vccd1
+ vccd1 _1377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4428_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[25\]
+ _0411_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\]
+ sky130_fd_sc_hd__dfstp_1
X_2689_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] _1336_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__a21boi_1
XANTENNA__2136__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4359_ clknet_leaf_11_wb_clk_i _0002_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4056__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_169_Left_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_178_Left_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2914__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_187_Left_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3630__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1991_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] net148 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__o22a_1
X_3730_ net246 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3661_ net269 vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload22 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_8
X_2612_ net195 _0909_ _1292_ _1290_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a32o_1
Xclkload11 clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__bufinv_16
X_3592_ net260 vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2543_ _0819_ team_10_WB.instance_to_wrap.host_col\[0\] _0851_ vssd1 vssd1 vccd1
+ vccd1 _1237_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_171_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4618__389 vssd1 vssd1 vccd1 vccd1 _4618__389/HI net389 sky130_fd_sc_hd__conb_1
X_2474_ net723 net129 _1211_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__o21a_1
X_4213_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[75\]
+ _0202_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[75\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4079__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4144_ clknet_leaf_28_wb_clk_i _0615_ _0143_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4075_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[6\]
+ _0095_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3026_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _1507_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[49\] sky130_fd_sc_hd__mux2_1
XANTENNA__3094__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3397__A2 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1995__A team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3928_ net268 vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload5 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_12
X_3859_ net269 vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout220 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] vssd1 vssd1 vccd1
+ vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout231 _0821_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_4
Xfanout242 net244 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_4
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
Xfanout253 net265 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_4
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_144_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout286 net289 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_4
Xfanout275 net285 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3388__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3625__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4221__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2190_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__or2_1
XANTENNA__4371__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1974_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\]
+ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__o22a_1
XANTENNA__3379__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4624__393 vssd1 vssd1 vccd1 vccd1 _4624__393/HI net393 sky130_fd_sc_hd__conb_1
XANTENNA__2423__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3713_ net250 vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3644_ net291 vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3000__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3575_ net282 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2526_ net520 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1
+ vccd1 vccd1 _0519_ sky130_fd_sc_hd__a22o_1
X_2457_ net549 net129 _1201_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o21a_1
Xhold17 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1
+ net473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold28 team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] vssd1 vssd1 vccd1 vccd1 net484
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ net5 net635 _1158_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__mux2_1
Xhold39 team_10_WB.instance_to_wrap.message_reg.msg\[6\] vssd1 vssd1 vccd1 vccd1 net495
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4127_ clknet_leaf_19_wb_clk_i _0598_ _0126_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_4058_ clknet_leaf_15_wb_clk_i _0543_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3009_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] net189 vssd1 vssd1 vccd1
+ vccd1 _1499_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4244__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4394__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2033__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3360_ team_10_WB.instance_to_wrap.host_row2\[57\] net180 net168 team_10_WB.instance_to_wrap.host_row2\[73\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2311_ _0841_ _1069_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__or3b_2
X_3291_ net295 _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__nor2_1
X_2242_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2173_ _0959_ _0962_ _0963_ _0937_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4117__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2272__A2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4267__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1957_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] net150 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__o22a_1
X_4676_ net182 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
X_1888_ net219 vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__inv_2
X_3627_ net248 vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3558_ net242 vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__inv_2
X_2509_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] net223 _1225_ vssd1
+ vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__and3_1
X_3489_ net253 vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
XANTENNA__2263__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4640__408 vssd1 vssd1 vccd1 vccd1 _4640__408/HI net408 sky130_fd_sc_hd__conb_1
XFILLER_0_66_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2860_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] _1450_ _1440_
+ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2791_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4530_ net341 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4461_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[18\]
+ _0444_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_159_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3412_ team_10_WB.instance_to_wrap.host_row1\[60\] _1704_ _1708_ team_10_WB.instance_to_wrap.host_row1\[76\]
+ _1787_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_123_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4392_ clknet_leaf_2_wb_clk_i _0777_ _0375_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_3343_ team_10_WB.instance_to_wrap.dispFSM.guesses\[24\] net171 _1704_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ net231 vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3274_ net534 _1660_ _1662_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_183_Right_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2225_ _0808_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__or3b_1
XANTENNA__2493__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2156_ _0949_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2087_ team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] net109 net135 net650 vssd1
+ vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2245__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2989_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\] net164 _1491_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[27\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_141_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4659_ net427 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4557__368 vssd1 vssd1 vccd1 vccd1 _4557__368/HI net368 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_150_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4432__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2236__A2 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4501__312 vssd1 vssd1 vccd1 vccd1 _4501__312/HI net312 sky130_fd_sc_hd__conb_1
XFILLER_0_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2010_ net219 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] net221 net222
+ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_29_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_X clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3961_ clknet_leaf_22_wb_clk_i _0481_ _0029_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_161_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2912_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\] net153 net121 net630
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[17\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3892_ net275 vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
X_2843_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] net475 net176
+ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2774_ net565 _1386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[27\]
+ sky130_fd_sc_hd__xor2_1
X_4513_ net324 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_170_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2935__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4305__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 net581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 net570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 team_10_WB.instance_to_wrap.dispFSM.guesses\[37\] vssd1 vssd1 vccd1 vccd1
+ net559 sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[1\]
+ _0427_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\]
+ sky130_fd_sc_hd__dfstp_1
Xhold147 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\] vssd1 vssd1 vccd1
+ vccd1 net603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 net69 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 team_10_WB.instance_to_wrap.dispFSM.guesses\[77\] vssd1 vssd1 vccd1 vccd1
+ net614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload21_A clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4375_ clknet_leaf_4_wb_clk_i _0760_ _0358_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[12\]
+ sky130_fd_sc_hd__dfstp_1
Xhold169 team_10_WB.instance_to_wrap.host_row1\[68\] vssd1 vssd1 vccd1 vccd1 net625
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3360__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3326_ team_10_WB.instance_to_wrap.host_row2\[80\] net173 net170 team_10_WB.instance_to_wrap.host_row2\[48\]
+ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__a221o_1
XANTENNA__3543__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4455__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3257_ _1651_ _1652_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout284_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ net297 net178 _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__nor3_2
XANTENNA__2466__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2208_ _0946_ net185 _0990_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__o21a_1
X_2139_ net134 _0934_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3103__A0 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2457__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4646__414 vssd1 vssd1 vccd1 vccd1 _4646__414/HI net414 sky130_fd_sc_hd__conb_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3406__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3972__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1968__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4328__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3628__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2490_ net511 net132 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] vssd1
+ vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4478__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3342__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4160_ clknet_leaf_30_wb_clk_i _0629_ _0149_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3111_ net535 net221 _1548_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4091_ clknet_leaf_12_wb_clk_i _0562_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3042_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] _1515_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[57\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3944_ clknet_leaf_3_wb_clk_i _0476_ net229 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3875_ net253 vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2826_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2757_ _1375_ _1376_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[20\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2688_ _1336_ _1337_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4427_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[24\]
+ _0410_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4358_ clknet_leaf_12_wb_clk_i _0001_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_input4_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _0815_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1679_ vssd1 vssd1
+ vccd1 vccd1 _1690_ sky130_fd_sc_hd__and3_1
X_4289_ clknet_leaf_18_wb_clk_i _0679_ _0278_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[12\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2439__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3100__A3 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3995__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3911__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1990_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] net149 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__o22a_1
XANTENNA__4150__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3660_ net294 vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload23 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__3012__C1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2611_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ _1291_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__or3_1
Xclkload12 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/X sky130_fd_sc_hd__clkbuf_8
X_3591_ net276 vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__inv_2
X_2542_ net225 _1068_ _1179_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__mux2_1
XANTENNA__2366__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4212_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[74\]
+ _0201_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[74\] sky130_fd_sc_hd__dfrtp_1
X_2473_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] net197 _1185_
+ _1210_ net130 vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__a221o_1
XFILLER_0_167_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4143_ clknet_leaf_9_wb_clk_i _0614_ _0142_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4074_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[5\]
+ _0094_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3025_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3032__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2054__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3927_ net289 vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3858_ net274 vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__inv_2
Xclkload6 clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_6
X_2809_ net230 _1414_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__nand2_1
X_3789_ net262 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout210 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\] vssd1 vssd1 vccd1
+ vccd1 net210 sky130_fd_sc_hd__buf_1
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_4
Xfanout221 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1 vccd1
+ vccd1 net221 sky130_fd_sc_hd__buf_2
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_4
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
Xfanout287 net289 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_4
Xfanout276 net280 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_4
Xfanout298 net7 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4173__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2899__A2 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2520__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2257__A team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1973_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0874_ _0879_ net159 vssd1
+ vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__o211a_1
X_3712_ net271 vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3643_ net288 vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4046__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3000__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3574_ net274 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3027__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2525_ net489 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1
+ vccd1 vccd1 _0520_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2456_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] net197 team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\]
+ net128 net130 vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__a221o_1
Xhold29 _0508_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 team_10_WB.instance_to_wrap.message_reg.msg\[5\] vssd1 vssd1 vccd1 vccd1 net474
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4196__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2387_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0856_ vssd1 vssd1 vccd1
+ vccd1 _1158_ sky130_fd_sc_hd__nand2_4
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4126_ clknet_leaf_20_wb_clk_i _0597_ _0125_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_4057_ clknet_leaf_15_wb_clk_i _0542_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3008_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\] net186 _1498_ net206
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[40\] sky130_fd_sc_hd__o211a_1
XANTENNA__3472__C1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout152_X net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3994__Q team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_X clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3290_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] _1668_ vssd1 vssd1 vccd1 vccd1
+ _1674_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2310_ team_10_WB.instance_to_wrap.host_col\[0\] _0859_ _0864_ vssd1 vssd1 vccd1
+ vccd1 _1086_ sky130_fd_sc_hd__or3b_1
XFILLER_0_57_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2241_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] _1022_ _1013_ _1015_
+ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__or4b_1
X_2172_ _0959_ _0962_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1956_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0874_ _0876_ net158 vssd1
+ vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4675_ net432 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1887_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 _0811_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout112_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3626_ net247 vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__inv_2
XANTENNA__2980__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3557_ net240 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
X_2508_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] _1224_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__o21a_2
X_3488_ net251 vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
X_2439_ net615 net133 _1191_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__a221o_1
X_4109_ clknet_leaf_9_wb_clk_i _0580_ _0108_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4211__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4361__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input42_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2487__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__C1 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2254__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2790_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4460_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[17\]
+ _0443_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2270__A team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2962__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3411_ team_10_WB.instance_to_wrap.host_row2\[52\] net171 _1784_ _1786_ vssd1 vssd1
+ vccd1 vccd1 _1787_ sky130_fd_sc_hd__a211o_1
X_4391_ clknet_leaf_5_wb_clk_i _0776_ _0374_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3342_ team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] net175 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[8\]
+ _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3273_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ vssd1 vssd1 vccd1 vccd1
+ _1663_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2224_ team_10_WB.EN_VAL_REG net41 _1008_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _0935_ _0948_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__or2_1
XFILLER_0_177_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2086_ team_10_WB.instance_to_wrap.dispFSM.guesses\[26\] net109 net136 net637 vssd1
+ vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4234__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4384__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2988_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\] net165 _1491_ net215
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[26\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1939_ team_10_WB.instance_to_wrap.host_message_reg.Cstate team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] _0861_ vssd1 vssd1 vccd1 vccd1
+ _0862_ sky130_fd_sc_hd__or4_2
X_4658_ net426 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__2953__A1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3609_ net276 vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4589_ net452 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2469__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4568__443 vssd1 vssd1 vccd1 vccd1 net443 _4568__443/LO sky130_fd_sc_hd__conb_1
XFILLER_0_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3433__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4540__351 vssd1 vssd1 vccd1 vccd1 _4540__351/HI net351 sky130_fd_sc_hd__conb_1
XFILLER_0_191_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4107__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3960_ clknet_leaf_23_wb_clk_i _0480_ _0028_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_161_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2911_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\] net155 net123 net710
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[16\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3424__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3891_ net281 vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2842_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] net176 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[0\] sky130_fd_sc_hd__and2b_1
XFILLER_0_170_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2773_ _1385_ _1386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[26\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4512_ net323 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XANTENNA__2935__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold126 team_10_WB.instance_to_wrap.host_row1\[42\] vssd1 vssd1 vccd1 vccd1 net582
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] vssd1 vssd1 vccd1
+ vccd1 net571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _0704_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold137 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net593 sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[0\]
+ _0426_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xhold148 team_10_WB.instance_to_wrap.host_row1\[78\] vssd1 vssd1 vccd1 vccd1 net604
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 team_10_WB.instance_to_wrap.host_row1\[74\] vssd1 vssd1 vccd1 vccd1 net615
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4374_ clknet_leaf_9_wb_clk_i _0759_ _0357_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3325_ team_10_WB.instance_to_wrap.host_row1\[64\] _1703_ net169 team_10_WB.instance_to_wrap.host_row1\[56\]
+ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__a22o_1
X_3256_ _0813_ _1650_ net295 vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2207_ net194 _0993_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__or2_1
XANTENNA__3112__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _0814_ _1607_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__or3b_4
XANTENNA_fanout277_A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2138_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ _0926_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__mux2_1
X_2069_ team_10_WB.instance_to_wrap.dispFSM.guesses\[43\] net112 net138 net636 vssd1
+ vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__o22a_1
XFILLER_0_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3415__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4524__335 vssd1 vssd1 vccd1 vccd1 _4524__335/HI net335 sky130_fd_sc_hd__conb_1
XFILLER_0_146_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1977__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3103__A1 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4611__385 vssd1 vssd1 vccd1 vccd1 _4611__385/HI net385 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_106_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3909__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1968__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3363__B _1740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ net553 net222 _1548_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__mux2_1
X_4090_ clknet_leaf_12_wb_clk_i _0561_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3041_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4508__319 vssd1 vssd1 vccd1 vccd1 _4508__319/HI net319 sky130_fd_sc_hd__conb_1
XFILLER_0_175_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3943_ net271 vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1959__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3874_ net252 vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__inv_2
X_2825_ net230 _1412_ _1417_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3030__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2756_ team_10_WB.instance_to_wrap.clock_div.count\[19\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ _1372_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2687_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] _1334_ _1319_ vssd1
+ vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4422__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4426_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[23\]
+ _0409_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_187_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2315__C_N net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4357_ clknet_leaf_11_wb_clk_i _0000_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3308_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net209 _1686_ _1688_
+ _1685_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__a41o_1
X_4288_ clknet_leaf_16_wb_clk_i _0678_ _0277_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_3239_ _1642_ _1611_ _1641_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__and3b_1
XANTENNA__3997__Q team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4445__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2262__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload24 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__clkinv_1
XTAP_TAPCELL_ROW_11_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload13 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_12
X_2610_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__or2_1
X_3590_ net252 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__inv_2
X_2541_ net224 _1236_ _1179_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__mux2_1
X_2472_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] net185 vssd1 vssd1 vccd1
+ vccd1 _1210_ sky130_fd_sc_hd__or2_1
X_4211_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[73\]
+ _0200_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[73\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3093__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4142_ clknet_leaf_20_wb_clk_i _0613_ _0141_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4073_ clknet_leaf_24_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[4\]
+ _0093_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3024_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] _1506_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[48\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_13_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3094__A3 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3926_ net286 vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_178_Right_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3857_ net273 vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload7 clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__clkinv_8
X_2808_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[2\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3788_ net293 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2739_ _1363_ _1364_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4409_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[6\]
+ _0392_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_1
Xfanout222 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\] vssd1 vssd1 vccd1
+ vccd1 net222 sky130_fd_sc_hd__buf_2
Xfanout211 team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1
+ net211 sky130_fd_sc_hd__buf_4
XANTENNA__3962__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_4
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout244 net266 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
Xfanout255 net258 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_4
Xfanout288 net289 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_4
Xfanout277 net280 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_4
Xfanout299 net300 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_2
Xfanout266 net298 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4318__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4468__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_21_wb_clk_i_X clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3481__X _1854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2257__B team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2036__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1972_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] net146 vssd1 vssd1 vccd1
+ vccd1 _0879_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_173_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4691_ net182 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
X_3711_ net236 vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3642_ net259 vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3985__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3573_ net281 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2524_ net494 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1
+ vccd1 vccd1 _0521_ sky130_fd_sc_hd__a22o_1
X_2455_ net507 net133 _1185_ _1200_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a22o_1
Xhold19 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\] vssd1 vssd1 vccd1
+ vccd1 net475 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] _1084_ _1156_
+ _1157_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__o22a_1
X_4125_ clknet_leaf_20_wb_clk_i _0596_ _0124_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3043__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4631__399 vssd1 vssd1 vccd1 vccd1 _4631__399/HI net399 sky130_fd_sc_hd__conb_1
X_4056_ clknet_leaf_15_wb_clk_i _0541_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3007_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] net190 vssd1 vssd1 vccd1
+ vccd1 _1498_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4171__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3909_ net248 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4140__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4290__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3917__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3652__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2240_ _1016_ _1017_ _1019_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__or4b_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2171_ team_10_WB.instance_to_wrap.correct\[2\] team_10_WB.instance_to_wrap.gamelogic.rights\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3454__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1955_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] net146 vssd1 vssd1 vccd1
+ vccd1 _0876_ sky130_fd_sc_hd__or2_1
XANTENNA__4013__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4674_ net183 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1886_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 _0810_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2450__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4163__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3625_ net248 vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__inv_2
X_3556_ net235 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__inv_2
X_2507_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] _1223_ vssd1 vssd1
+ vccd1 vccd1 _1224_ sky130_fd_sc_hd__or2_1
X_3487_ net267 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2438_ net579 net133 _1191_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__a221o_1
X_2369_ _0871_ _1143_ _1087_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__a21oi_1
X_4108_ clknet_leaf_11_wb_clk_i _0579_ _0107_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_4039_ clknet_leaf_22_wb_clk_i _0524_ _0080_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2248__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1931__B1 team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input35_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3436__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2239__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1998__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4036__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4186__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2270__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2962__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4390_ clknet_leaf_4_wb_clk_i _0775_ _0373_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[27\]
+ sky130_fd_sc_hd__dfstp_1
X_3410_ team_10_WB.instance_to_wrap.host_row1\[68\] _1703_ net180 team_10_WB.instance_to_wrap.host_row2\[60\]
+ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__a221o_1
X_3341_ team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] net173 net181 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\]
+ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3272_ net295 _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2223_ net42 net40 net43 _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _0822_ net217 _0948_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2085_ team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] net112 net139 net683 vssd1
+ vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__o22a_1
XFILLER_0_177_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2445__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_wb_clk_i_X clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_158_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1989__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2987_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] net165 _1491_ net216
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[25\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3557__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1938_ _0840_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__nand2_1
X_4657_ net425 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_140_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1869_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] vssd1 vssd1 vccd1 vccd1
+ _0794_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3608_ net281 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4588_ net451 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_149_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3539_ net246 vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__inv_2
XANTENNA__4059__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3418__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2636__A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_73_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input38_X net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3409__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2910_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\] net157 _1472_ net594
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[15\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3890_ net274 vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2841_ _1010_ _1238_ _1241_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2772_ team_10_WB.instance_to_wrap.clock_div.count\[25\] team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ team_10_WB.instance_to_wrap.clock_div.count\[26\] _1382_ vssd1 vssd1 vccd1 vccd1
+ _1386_ sky130_fd_sc_hd__and4_1
X_4511_ net322 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_170_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2935__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4442_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[39\]
+ _0425_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold116 team_10_WB.instance_to_wrap.host_row1\[69\] vssd1 vssd1 vccd1 vccd1 net572
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_91_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold105 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 net561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold138 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\] vssd1 vssd1 vccd1
+ vccd1 net594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] vssd1 vssd1 vccd1 vccd1
+ net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 team_10_WB.instance_to_wrap.dispFSM.guesses\[21\] vssd1 vssd1 vccd1 vccd1
+ net583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4373_ clknet_leaf_2_wb_clk_i _0758_ _0356_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3360__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3324_ _1681_ _1698_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__and2_2
XFILLER_0_21_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3255_ _0813_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__nor2_1
XANTENNA__4201__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2206_ net194 _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_185_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\]
+ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__and3_1
XANTENNA__3051__S net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2137_ net134 _0933_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__and2_1
XANTENNA__4351__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2068_ team_10_WB.instance_to_wrap.dispFSM.guesses\[44\] net112 net138 net687 vssd1
+ vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4563__374 vssd1 vssd1 vccd1 vccd1 _4563__374/HI net374 sky130_fd_sc_hd__conb_1
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3351__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4581__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4224__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3660__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4374__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] _1514_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[56\] sky130_fd_sc_hd__mux2_1
XFILLER_0_65_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4547__358 vssd1 vssd1 vccd1 vccd1 _4547__358/HI net358 sky130_fd_sc_hd__conb_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ net251 vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3873_ net252 vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2824_ _1418_ _1426_ _1407_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_14_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_143_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2755_ team_10_WB.instance_to_wrap.clock_div.count\[20\] _1374_ vssd1 vssd1 vccd1
+ vccd1 _1375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2686_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\]
+ _1332_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4425_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[22\]
+ _0408_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3333__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4356_ clknet_leaf_22_wb_clk_i _0746_ _0345_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_3307_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_6_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4287_ clknet_leaf_22_wb_clk_i _0677_ _0276_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3570__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3238_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ _1638_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__and3_1
X_3169_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1551_ _1595_ vssd1 vssd1 vccd1
+ vccd1 _0500_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_138_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_11_wb_clk_i_X clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4247__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4397__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4652__420 vssd1 vssd1 vccd1 vccd1 _4652__420/HI net420 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_147_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4576__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_156_Left_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2543__B team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_184_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload25 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_8
Xclkload14 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_11_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2540_ _0818_ _0842_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__nor2_1
X_2471_ net518 net129 _1194_ _1209_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__o22a_1
X_4210_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[72\]
+ _0199_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[72\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4141_ clknet_leaf_11_wb_clk_i _0612_ _0140_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4072_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[3\]
+ _0092_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3023_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3925_ net255 vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__inv_2
XANTENNA__2054__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3856_ net274 vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__inv_2
Xclkload8 clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_8
X_2807_ _1413_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__inv_2
XANTENNA__3003__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3787_ net261 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout302_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2738_ team_10_WB.instance_to_wrap.clock_div.count\[13\] team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ _1362_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4636__404 vssd1 vssd1 vccd1 vccd1 _4636__404/HI net404 sky130_fd_sc_hd__conb_1
X_4408_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[5\]
+ _0391_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2669_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] _1321_ _1319_ vssd1
+ vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__o21ai_1
Xfanout201 net63 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout223 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\] vssd1 vssd1 vccd1
+ vccd1 net223 sky130_fd_sc_hd__clkbuf_2
Xfanout212 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1
+ net212 sky130_fd_sc_hd__buf_4
X_4339_ clknet_leaf_15_wb_clk_i _0729_ _0328_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[62\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout234 net266 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
Xfanout245 net249 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_4
Xfanout256 net258 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_4
XFILLER_0_157_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_4
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_4
Xfanout267 net275 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_4
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4412__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1971_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] net148 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3710_ net236 vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__inv_2
X_4690_ net437 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_173_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ net287 vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__inv_2
X_3572_ net288 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2523_ net493 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1
+ vccd1 vccd1 _0522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2454_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] net186 vssd1 vssd1 vccd1
+ vccd1 _1200_ sky130_fd_sc_hd__or2_1
X_2385_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__a21o_1
X_4124_ clknet_leaf_20_wb_clk_i _0595_ _0123_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput1 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
X_4055_ clknet_leaf_15_wb_clk_i _0540_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_143_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4092__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3006_ net211 net126 _1496_ net735 net160 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[39\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout252_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3908_ net290 vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3839_ net287 vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4435__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3189__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3933__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2170_ _0961_ _0960_ _0959_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4665__430 vssd1 vssd1 vccd1 vccd1 _4665__430/HI net430 sky130_fd_sc_hd__conb_1
XFILLER_0_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3952__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4272__Q team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_1954_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4673_ net182 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1885_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 _0809_ sky130_fd_sc_hd__inv_2
X_3624_ net248 vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__inv_2
XANTENNA__4308__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2193__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3555_ net235 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__inv_2
X_3486_ _1409_ _1436_ _1438_ _1405_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__o211a_1
XANTENNA__3390__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2506_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__or4_1
X_2437_ net519 net133 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__a22o_1
XANTENNA__4458__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2368_ _1091_ _1137_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__xor2_1
X_4107_ clknet_leaf_10_wb_clk_i _0578_ _0106_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2299_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__inv_2
XANTENNA__3445__A1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4038_ clknet_leaf_21_wb_clk_i _0523_ _0079_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2487__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3436__A1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2239__A2 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3975__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1998__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1998__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3340_ _1694_ _1718_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__nor2_4
XANTENNA__3372__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4591__454 vssd1 vssd1 vccd1 vccd1 net454 _4591__454/LO sky130_fd_sc_hd__conb_1
XFILLER_0_110_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ vssd1 vssd1 vccd1 vccd1
+ _1661_ sky130_fd_sc_hd__and4_1
X_2222_ net182 vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__inv_2
XANTENNA__2478__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2084_ team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] net112 net139 net649 vssd1
+ vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4130__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2938__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2986_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] net164 _1491_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[24\]
+ sky130_fd_sc_hd__o22a_1
X_1937_ _0842_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__nor2_1
X_4656_ net424 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_138_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1868_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1 vccd1 vccd1
+ _0793_ sky130_fd_sc_hd__inv_2
X_4587_ net201 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_3607_ net282 vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__inv_2
XANTENNA__4280__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3538_ net246 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2189__A team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3469_ team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] net180 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[71\]
+ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3998__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_191_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3354__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4003__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4153__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2840_ _1405_ _1426_ _1437_ _1410_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2771_ team_10_WB.instance_to_wrap.clock_div.count\[26\] _1384_ vssd1 vssd1 vccd1
+ vccd1 _1385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4510_ net321 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4441_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[38\]
+ _0424_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\] vssd1 vssd1 vccd1
+ vccd1 net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 team_10_WB.instance_to_wrap.dispFSM.guesses\[45\] vssd1 vssd1 vccd1 vccd1
+ net573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold139 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[15\] vssd1 vssd1
+ vccd1 vccd1 net595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\] vssd1 vssd1 vccd1 vccd1
+ net584 sky130_fd_sc_hd__dlygate4sd3_1
X_4372_ clknet_leaf_7_wb_clk_i _0757_ _0355_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ sky130_fd_sc_hd__dfstp_2
X_3323_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ _1698_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__and3_2
XFILLER_0_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3254_ net632 _1609_ _1650_ net230 vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2205_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] vssd1 vssd1 vccd1 vccd1 _0993_
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_185_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _1608_
+ sky130_fd_sc_hd__and3_1
X_2136_ net216 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0933_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout165_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2067_ net739 net143 net108 net573 vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2191__B team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2969_ team_10_WB.instance_to_wrap.gamelogic.letter\[7\] net126 _1482_ net617 net160
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[15\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3336__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4639_ net407 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2066__B1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3941_ net254 vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3872_ net252 vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__inv_2
X_2823_ _0514_ _0513_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2754_ _1373_ _1374_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[19\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4049__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2685_ _1334_ _1335_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[8\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4424_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[21\]
+ _0407_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_4355_ clknet_leaf_16_wb_clk_i _0745_ _0344_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[78\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4199__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3306_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__nand2b_2
XANTENNA__3851__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4286_ clknet_leaf_18_wb_clk_i _0676_ _0275_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_3237_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ _1637_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] vssd1 vssd1 vccd1 vccd1
+ _1641_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_146_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3062__S net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4530__341 vssd1 vssd1 vccd1 vccd1 _4530__341/HI net341 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3168_ _1586_ _1590_ _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__a21o_1
XFILLER_0_178_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2119_ _0920_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_65_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3099_ _0789_ net206 vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout168_X net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3254__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_X clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload26 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__3012__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload15 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_11_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4341__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2470_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] net197 team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ net126 vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_192_Right_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4140_ clknet_leaf_11_wb_clk_i _0611_ _0139_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2523__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4514__325 vssd1 vssd1 vccd1 vccd1 _4514__325/HI net325 sky130_fd_sc_hd__conb_1
XANTENNA__4491__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4071_ clknet_leaf_24_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[2\]
+ _0091_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3022_ net541 net185 _1505_ net202 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[47\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_182_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3484__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4275__Q team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3924_ net290 vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3855_ net273 vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload9 clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_12
XFILLER_0_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2806_ net230 _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__nand2_1
X_3786_ net280 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__inv_2
X_4601__375 vssd1 vssd1 vccd1 vccd1 _4601__375/HI net375 sky130_fd_sc_hd__conb_1
X_4675__432 vssd1 vssd1 vccd1 vccd1 _4675__432/HI net432 sky130_fd_sc_hd__conb_1
X_2737_ team_10_WB.instance_to_wrap.clock_div.count\[13\] _1362_ net725 vssd1 vssd1
+ vccd1 vccd1 _1363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2668_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] _1321_ vssd1 vssd1
+ vccd1 vccd1 _1324_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4407_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[4\]
+ _0390_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2599_ _0903_ _1280_ _1282_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__and3b_1
Xfanout213 team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1
+ net213 sky130_fd_sc_hd__buf_4
Xfanout202 net203 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_4
Xfanout224 team_10_WB.instance_to_wrap.host_col\[2\] vssd1 vssd1 vccd1 vccd1 net224
+ sky130_fd_sc_hd__clkbuf_2
Xfanout246 net249 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_4
X_4338_ clknet_leaf_20_wb_clk_i _0728_ _0327_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout268 net275 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
Xfanout279 net280 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_4
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
XFILLER_0_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4269_ clknet_leaf_0_wb_clk_i _0659_ _0258_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_2_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4214__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4364__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4587__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3491__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1970_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] net149 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2441__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2992__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4659__427 vssd1 vssd1 vccd1 vccd1 _4659__427/HI net427 sky130_fd_sc_hd__conb_1
X_3640_ net259 vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__inv_2
X_3571_ net242 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__inv_2
X_2522_ net486 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1
+ vccd1 vccd1 _0523_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2453_ net554 net133 _1185_ _1199_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__a22o_1
X_2384_ _1154_ _1155_ _1087_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__a21oi_1
X_4123_ clknet_leaf_28_wb_clk_i _0594_ _0122_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_4054_ clknet_leaf_15_wb_clk_i _0539_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput2 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_143_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3005_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\] net164 _1497_ net212
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[38\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3472__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4387__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout245_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3907_ net255 vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__inv_2
X_3838_ net286 vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_175_Left_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3769_ net284 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__inv_2
XANTENNA__2196__C1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2499__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_184_Left_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3463__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3311__A_N net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_193_Left_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2974__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3151__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3454__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1953_ net147 net159 vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__nand2_2
XFILLER_0_189_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4672_ net182 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1884_ team_10_WB.instance_to_wrap.message_reg.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _0808_ sky130_fd_sc_hd__inv_2
XANTENNA__2965__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3623_ net237 vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3554_ net235 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__inv_2
X_2505_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[1\] vssd1 vssd1 vccd1 vccd1 _1222_
+ sky130_fd_sc_hd__and3b_1
X_3485_ net538 _1284_ net195 vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__o21a_1
X_2436_ _1193_ _1194_ net527 net131 vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2367_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] _1084_ _1140_
+ _1142_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__o22a_1
X_4106_ clknet_leaf_11_wb_clk_i _0577_ _0105_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_2298_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _0823_ _1069_ vssd1 vssd1
+ vccd1 vccd1 _1077_ sky130_fd_sc_hd__nand3_2
X_4037_ clknet_leaf_22_wb_clk_i _0522_ _0078_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout150_X net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4607__381 vssd1 vssd1 vccd1 vccd1 _4607__381/HI net381 sky130_fd_sc_hd__conb_1
XFILLER_0_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4402__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3381__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__A2 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1998__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4082__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3270_ net295 _1659_ _1660_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__nor3_1
XFILLER_0_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _1001_ _1002_ _1003_ _1006_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__or4_1
X_2152_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2083_ net559 net143 net108 net605 vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1989__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2938__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2985_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1936_ net228 _0857_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__or3b_2
XFILLER_0_56_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1867_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] vssd1 vssd1 vccd1 vccd1
+ _0792_ sky130_fd_sc_hd__inv_2
XANTENNA__4425__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4655_ net423 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA_fanout208_A team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3606_ net281 vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout110_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4586_ net199 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3537_ net246 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3468_ net464 net177 _1841_ net229 vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__o211a_1
XANTENNA__2189__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3115__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3399_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] _1688_ _1679_ net209
+ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2419_ net203 _0942_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_30_wb_clk_i_X clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2636__C _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3051__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input40_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4368__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4595__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3409__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4448__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3042__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ _1383_ _1384_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[25\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4440_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[37\]
+ _0423_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold107 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 net563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold118 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\] vssd1 vssd1 vccd1
+ vccd1 net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 team_10_WB.instance_to_wrap.dispFSM.guesses\[79\] vssd1 vssd1 vccd1 vccd1
+ net585 sky130_fd_sc_hd__dlygate4sd3_1
X_4371_ clknet_leaf_9_wb_clk_i _0756_ _0354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_21_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3322_ _1683_ _1694_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3253_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] _1607_ _1609_ vssd1 vssd1
+ vccd1 vccd1 _1650_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3184_ _1603_ _1604_ _1605_ _1606_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__or4_1
X_2204_ _0946_ net194 _0990_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_185_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ net134 _0932_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2066_ team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] net114 net142 net717 vssd1
+ vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout158_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2472__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2968_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] net165 _1483_ net212
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[14\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1919_ net224 net225 team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1
+ vccd1 _0842_ sky130_fd_sc_hd__or3_2
X_4638_ net406 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
X_2899_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\] net152 net124 net591
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[4\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ net444 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_12_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3024__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4120__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4270__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3940_ net290 vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4627__395 vssd1 vssd1 vccd1 vccd1 _4627__395/HI net395 sky130_fd_sc_hd__conb_1
X_3871_ net253 vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_176_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2822_ net296 _1417_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2753_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[19\]
+ team_10_WB.instance_to_wrap.clock_div.count\[18\] _1367_ vssd1 vssd1 vccd1 vccd1
+ _1374_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_14_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3988__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2684_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] _1332_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4423_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[20\]
+ _0406_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_4354_ clknet_leaf_20_wb_clk_i _0744_ _0343_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_3305_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__and2b_2
XANTENNA_clkload12_A clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4285_ clknet_leaf_16_wb_clk_i _0675_ _0274_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_3236_ net610 _1638_ _1640_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_146_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout275_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3167_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1278_ _1568_ _1593_ vssd1 vssd1
+ vccd1 vccd1 _1594_ sky130_fd_sc_hd__a211o_1
XFILLER_0_178_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2118_ team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] team_10_WB.instance_to_wrap.buffer.temp_guess\[6\]
+ team_10_WB.instance_to_wrap.buffer.temp_guess\[5\] team_10_WB.instance_to_wrap.buffer.temp_guess\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__or4_1
X_3098_ net197 net743 net185 _1543_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[85\]
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_166_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ net597 net144 net107 net624 vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4143__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4293__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3088__A3 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/X sky130_fd_sc_hd__clkbuf_8
Xclkload27 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_11_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4553__364 vssd1 vssd1 vccd1 vccd1 _4553__364/HI net364 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_79_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4070_ clknet_leaf_24_wb_clk_i net476 _0090_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3021_ _0796_ net185 vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2039__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4016__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3923_ net254 vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3854_ net273 vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2805_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[1\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3785_ net284 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
XANTENNA__4166__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2736_ team_10_WB.instance_to_wrap.clock_div.count\[13\] _1362_ vssd1 vssd1 vccd1
+ vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[13\] sky130_fd_sc_hd__xor2_1
XFILLER_0_14_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2667_ _1318_ _1322_ _1323_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[2\]
+ sky130_fd_sc_hd__and3_1
X_4406_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[3\]
+ _0389_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_97_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2598_ _1275_ _1278_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__or2_1
Xfanout214 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1
+ net214 sky130_fd_sc_hd__clkbuf_4
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlymetal6s2s_1
X_4337_ clknet_leaf_19_wb_clk_i _0727_ _0326_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[60\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout236 net237 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_4
Xfanout225 team_10_WB.instance_to_wrap.host_col\[1\] vssd1 vssd1 vccd1 vccd1 net225
+ sky130_fd_sc_hd__buf_2
Xfanout247 net248 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_4
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_4
X_4268_ clknet_leaf_5_wb_clk_i _0658_ _0257_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout258 net265 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2197__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ net172 vssd1
+ vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout180_X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3475__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4199_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[61\]
+ _0188_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[61\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4496__307 vssd1 vssd1 vccd1 vccd1 _4496__307/HI net307 sky130_fd_sc_hd__conb_1
XFILLER_0_134_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4537__348 vssd1 vssd1 vccd1 vccd1 _4537__348/HI net348 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_170_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4039__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4189__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3570_ net240 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__inv_2
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2521_ net474 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] vssd1 vssd1
+ vccd1 vccd1 _0524_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1952__B1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2452_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] net186 vssd1 vssd1 vccd1
+ vccd1 _1199_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2383_ _1123_ _1127_ _1136_ _0871_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o31a_1
X_4122_ clknet_leaf_20_wb_clk_i _0593_ _0121_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_4053_ clknet_leaf_15_wb_clk_i _0538_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_143_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3004_ _1484_ _1496_ _1497_ _1493_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[37\]
+ sky130_fd_sc_hd__a22oi_1
Xinput3 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4642__410 vssd1 vssd1 vccd1 vccd1 _4642__410/HI net410 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_102_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3906_ net272 vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout238_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2480__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3837_ net247 vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3768_ net278 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2719_ _1351_ _1352_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3699_ net245 vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3448__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4331__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4481__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3384__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3007__A team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3439__A0 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1952_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0874_ net158 _0863_ vssd1
+ vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4671_ net183 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1883_ team_10_WB.instance_to_wrap.message_reg.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _0807_ sky130_fd_sc_hd__inv_2
XFILLER_0_189_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3622_ net244 vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_190_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4559__370 vssd1 vssd1 vccd1 vccd1 _4559__370/HI net370 sky130_fd_sc_hd__conb_1
X_3553_ net256 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__inv_2
X_3484_ net539 net177 _1856_ net229 vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2504_ net222 _1221_ _1217_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__mux2_1
XANTENNA__4204__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2435_ net131 _1190_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ clknet_leaf_9_wb_clk_i _0576_ _0104_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2366_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout188_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2297_ _1069_ _1074_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__or2_1
XANTENNA__4354__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_20_wb_clk_i_X clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4036_ clknet_leaf_22_wb_clk_i _0521_ _0077_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2653__B2 _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2503__A_N net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3372__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ net32 net31 _1004_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__or4_1
XANTENNA__4377__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2151_ net162 _0918_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2082_ team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] net114 net140 net724 vssd1
+ vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_49_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_187_Right_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2984_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] _1191_ _1489_ _1490_
+ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_32_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2938__A2 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1935_ _0847_ net196 vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__nand2_2
XFILLER_0_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4654_ net422 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_138_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1866_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1
+ _0791_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_15_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3605_ net291 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__inv_2
X_4585_ net200 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
X_3536_ net246 vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__inv_2
X_3467_ net169 _1839_ _1840_ _1838_ _1403_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_149_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3398_ team_10_WB.instance_to_wrap.host_row2\[43\] team_10_WB.instance_to_wrap.dispFSM.guesses\[19\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__mux2_1
X_2418_ _1178_ _1179_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_24_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2349_ _1122_ _1102_ _1117_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__and3b_1
X_4019_ clknet_leaf_29_wb_clk_i _0504_ _0066_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.unlocked
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3354__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input33_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4384__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_51_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold108 team_10_WB.instance_to_wrap.dispFSM.guesses\[61\] vssd1 vssd1 vccd1 vccd1
+ net564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\] vssd1 vssd1 vccd1
+ vccd1 net575 sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ clknet_leaf_29_wb_clk_i _0755_ _0353_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3321_ _1686_ _1695_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__and2_2
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_60_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3252_ _1610_ _1649_ net295 vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3183_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__or4bb_1
X_2203_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.correct\[0\]
+ team_10_WB.instance_to_wrap.correct\[2\] vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__and3b_1
XANTENNA__1922__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2134_ net215 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2065_ team_10_WB.instance_to_wrap.dispFSM.guesses\[55\] net143 net108 net568 vssd1
+ vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_16_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2967_ _1479_ _1483_ _1484_ _1482_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[13\]
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2898_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\] net153 net121 net603
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[3\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1918_ team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4637_ net405 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3336__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3076__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4568_ net443 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_12_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2544__A0 team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4499_ net310 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
X_3519_ net233 vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4072__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4379__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3015__A team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4415__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3870_ net253 vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2821_ _1405_ _1424_ _1425_ _1411_ _1419_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2752_ team_10_WB.instance_to_wrap.clock_div.count\[19\] _1372_ vssd1 vssd1 vccd1
+ vccd1 _1373_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2683_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] _1332_ vssd1 vssd1
+ vccd1 vccd1 _1334_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4422_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[19\]
+ _0405_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_4353_ clknet_leaf_18_wb_clk_i _0743_ _0342_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[76\]
+ sky130_fd_sc_hd__dfstp_1
X_3304_ _0815_ net209 _1679_ _1681_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__and4_1
X_4284_ clknet_leaf_19_wb_clk_i net483 _0273_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3235_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\] _1638_ _1612_ vssd1
+ vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_146_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4095__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3166_ _0891_ _0899_ _0906_ net227 vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2117_ team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] team_10_WB.instance_to_wrap.buffer.temp_guess\[2\]
+ team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__or4_1
X_3097_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] net203 vssd1 vssd1 vccd1
+ vccd1 _1543_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2048_ team_10_WB.instance_to_wrap.dispFSM.guesses\[64\] net115 net141 net676 vssd1
+ vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_105_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout268_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3006__B2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3006__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3999_ clknet_leaf_27_wb_clk_i net457 net254 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_107_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4438__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload17 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/X sky130_fd_sc_hd__clkbuf_8
Xclkload28 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_4
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3020_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\] net186 _1504_ net205
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[46\] sky130_fd_sc_hd__o211a_1
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2039__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3955__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3922_ net272 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3853_ net250 vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__inv_2
XFILLER_0_183_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2804_ _1405_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__nor2_1
XANTENNA__1928__A team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3784_ net279 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2735_ _1361_ _1362_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2666_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1323_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1970__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4405_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[2\]
+ _0388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_4336_ clknet_leaf_17_wb_clk_i _0726_ _0325_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[59\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2597_ _1275_ _1278_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__nor2_1
Xfanout204 team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 net204
+ sky130_fd_sc_hd__clkbuf_4
Xfanout237 net266 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_4
Xfanout226 _0897_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
Xfanout215 team_10_WB.instance_to_wrap.gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1
+ net215 sky130_fd_sc_hd__buf_4
X_4267_ clknet_leaf_5_wb_clk_i _0657_ _0256_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1950__X _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_4
Xfanout259 net261 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_4
X_3218_ net711 _1626_ _1629_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o21a_1
X_4198_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[60\]
+ _0187_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[60\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_31_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_2_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3149_ _0903_ _1277_ _1280_ _1578_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout173_X net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4110__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1961__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold280 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\] vssd1 vssd1 vccd1
+ vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3978__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4392__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3439__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4520__331 vssd1 vssd1 vccd1 vccd1 _4520__331/HI net331 sky130_fd_sc_hd__conb_1
XFILLER_0_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2520_ net495 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1
+ vccd1 vccd1 _0525_ sky130_fd_sc_hd__a22o_1
X_2451_ net551 net131 _1185_ _1198_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1952__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2382_ _1123_ _1136_ _1127_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__o21ai_1
X_4121_ clknet_leaf_20_wb_clk_i _0592_ _0120_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_4052_ clknet_leaf_15_wb_clk_i _0537_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_X clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_127_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3003_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\] net164 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[4\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[36\]
+ sky130_fd_sc_hd__o22a_1
Xinput4 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4133__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3905_ net287 vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3836_ net286 vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout133_A _1183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4283__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3767_ net278 vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3393__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2718_ net533 _1349_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3698_ net245 vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__inv_2
X_2649_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4319_ clknet_leaf_18_wb_clk_i _0709_ _0308_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_161_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4504__315 vssd1 vssd1 vccd1 vccd1 _4504__315/HI net315 sky130_fd_sc_hd__conb_1
XFILLER_0_107_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4387__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4006__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3007__B net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4156__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1951_ team_10_WB.instance_to_wrap.host_message_reg.Cstate team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] _0861_ vssd1 vssd1 vccd1 vccd1
+ _0874_ sky130_fd_sc_hd__nor4_4
X_1882_ team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
X_4670_ net182 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3621_ net237 vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3375__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3552_ net256 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2503_ net222 _0889_ net221 vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__and3b_1
XANTENNA__1925__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3483_ _1847_ _1853_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2434_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] _1192_ vssd1 vssd1 vccd1
+ vccd1 _1193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2365_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _0823_ _1069_ _1085_
+ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__a31o_1
X_4104_ clknet_leaf_25_wb_clk_i _0575_ _0103_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2296_ _0841_ _1069_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__or2_2
X_4035_ clknet_leaf_22_wb_clk_i _0520_ _0076_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3079__S net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3819_ net247 vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__inv_2
XANTENNA__3366__B1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4179__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4649__417 vssd1 vssd1 vccd1 vccd1 _4649__417/HI net417 sky130_fd_sc_hd__conb_1
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3357__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3018__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2150_ net162 _0918_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nor2_1
X_2081_ team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] net144 net107 net611 vssd1
+ vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2983_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\]
+ _0836_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net165 vssd1 vssd1 vccd1
+ vccd1 _1490_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_32_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1934_ _0843_ net196 vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4653_ net421 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
Xinput40 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
X_1865_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\] vssd1 vssd1 vccd1 vccd1
+ _0790_ sky130_fd_sc_hd__inv_2
XANTENNA__2531__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3604_ net291 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__inv_2
X_4584_ net199 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3535_ net246 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__inv_2
X_3466_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1686_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ net209 vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__and4b_1
XANTENNA__4321__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2417_ _1164_ _1167_ _1168_ _1169_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3397_ team_10_WB.instance_to_wrap.host_row1\[59\] _1704_ _1768_ _1773_ vssd1 vssd1
+ vccd1 vccd1 _1774_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2348_ _1102_ _1117_ _1122_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__and3b_1
XANTENNA__4471__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2279_ _0917_ _0948_ _1034_ _1047_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__o31ai_1
X_4018_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[2\]
+ net243 vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4620__391 vssd1 vssd1 vccd1 vccd1 _4620__391/HI net391 sky130_fd_sc_hd__conb_1
XFILLER_0_132_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input26_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4344__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold109 team_10_WB.instance_to_wrap.clock_div.count\[27\] vssd1 vssd1 vccd1 vccd1
+ net565 sky130_fd_sc_hd__dlygate4sd3_1
X_3320_ team_10_WB.instance_to_wrap.host_row2\[40\] net174 _1699_ team_10_WB.instance_to_wrap.host_row1\[48\]
+ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3251_ _1609_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_119_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3182_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 _1605_
+ sky130_fd_sc_hd__or3b_1
X_2202_ _0918_ _0972_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2133_ net134 _0931_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__and2_1
X_2064_ team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] net114 net140 net660 vssd1
+ vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2966_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] _1192_ vssd1 vssd1 vccd1
+ vccd1 _1484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2897_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\] net152 net124 net574
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[2\]
+ sky130_fd_sc_hd__o22a_1
X_1917_ team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout213_A team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4636_ net404 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_114_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4567_ net442 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4498_ net309 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
X_3518_ net232 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3449_ _1821_ _1822_ _1823_ net301 vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__o31a_1
XFILLER_0_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4685__436 vssd1 vssd1 vccd1 vccd1 _4685__436/HI net436 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_68_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4217__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4367__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2960__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3015__B net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2820_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2751_ _1371_ _1372_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[18\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2682_ _1318_ _1331_ _1333_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[7\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4421_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[18\]
+ _0404_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_96_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4352_ clknet_leaf_18_wb_clk_i _0742_ _0341_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[75\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2526__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4283_ clknet_leaf_15_wb_clk_i _0673_ _0272_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_3303_ _1680_ _1683_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__nor2_1
X_3234_ net526 _1637_ _1639_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_146_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3165_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] _1551_ _1591_ _1592_ vssd1 vssd1
+ vccd1 vccd1 _0499_ sky130_fd_sc_hd__o22a_1
X_3096_ net207 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] net191 _1542_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[84\] sky130_fd_sc_hd__a31o_1
X_2116_ net159 _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__or2_2
X_2047_ team_10_WB.instance_to_wrap.dispFSM.guesses\[65\] net109 net136 net662 vssd1
+ vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_65_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3006__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3998_ clknet_leaf_27_wb_clk_i net459 net254 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2949_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] net163 _1478_ net216 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[1\] sky130_fd_sc_hd__o22a_1
XFILLER_0_91_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1973__C1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2004__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4619_ net390 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_187_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2453__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3786__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload18 clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_6
Xclkload29 clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3313__X _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3484__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3921_ net286 vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__inv_2
XANTENNA__2444__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3852_ net289 vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2803_ _1407_ _0517_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_193_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3783_ net279 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2734_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] _1356_ vssd1 vssd1 vccd1 vccd1
+ _1362_ sky130_fd_sc_hd__and4_1
X_2665_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4404_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[1\]
+ _0387_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2596_ _1276_ _1280_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__nand2_1
XANTENNA__4062__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 net208 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_4
X_4335_ clknet_leaf_22_wb_clk_i _0725_ _0324_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[58\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout238 net240 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_4
Xfanout227 _0897_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_1
Xfanout216 team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1
+ net216 sky130_fd_sc_hd__buf_4
X_4266_ clknet_leaf_5_wb_clk_i _0656_ _0255_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout249 net265 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
XFILLER_0_66_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3217_ net172 _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__nor2_1
X_4197_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[59\]
+ _0186_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[59\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3475__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3148_ _1571_ _1577_ _1560_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__mux2_1
XANTENNA__3350__C_N net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3079_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout166_X net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2986__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4405__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1961__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold270 team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] vssd1 vssd1 vccd1 vccd1
+ net726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold281 team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] vssd1 vssd1 vccd1 vccd1
+ net737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2977__B2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2450_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\] net186 vssd1 vssd1 vccd1
+ vccd1 _1198_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_93_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2381_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] _1084_ _1141_
+ _1153_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__o22a_1
X_4120_ clknet_leaf_28_wb_clk_i net509 _0119_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_4051_ clknet_leaf_15_wb_clk_i _0536_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3457__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3002_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\] net163 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[35\]
+ sky130_fd_sc_hd__o22a_1
Xinput5 gpio_in[28] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_2
XFILLER_0_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_6_wb_clk_i_X clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3904_ net267 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__inv_2
XANTENNA__2968__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2534__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4428__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3835_ net247 vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__inv_2
X_3766_ net293 vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2717_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ team_10_WB.instance_to_wrap.clock_div.count\[6\] _1347_ vssd1 vssd1 vccd1 vccd1
+ _1351_ sky130_fd_sc_hd__and4_1
XANTENNA__3365__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3697_ net245 vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_144_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2648_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[1\] vssd1 vssd1 vccd1 vccd1 _1310_
+ sky130_fd_sc_hd__or3b_2
X_2579_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] _1259_ _0904_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_77_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4318_ clknet_leaf_19_wb_clk_i _0708_ _0307_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[41\]
+ sky130_fd_sc_hd__dfstp_1
X_4249_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[5\]
+ _0238_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3448__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_153_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3081__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4543__354 vssd1 vssd1 vccd1 vccd1 _4543__354/HI net354 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_172_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_162_Left_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3945__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input11_X net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_171_Left_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3072__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1950_ _0841_ _0871_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__or2_2
X_1881_ team_10_WB.instance_to_wrap.gamelogic.green vssd1 vssd1 vccd1 vccd1 _0806_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3620_ net241 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_180_Left_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3551_ net256 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__inv_2
X_2502_ net221 _1220_ _1217_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__mux2_1
XANTENNA__1925__A2 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3482_ net179 _1854_ _1403_ _1689_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2433_ net604 net132 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2364_ _1138_ _1139_ _1088_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__o21a_1
X_4103_ clknet_leaf_24_wb_clk_i _0574_ _0102_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2529__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4100__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2295_ _0840_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4034_ clknet_leaf_22_wb_clk_i _0519_ _0075_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2102__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4527__338 vssd1 vssd1 vccd1 vccd1 _4527__338/HI net338 sky130_fd_sc_hd__conb_1
XFILLER_0_176_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4250__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3818_ net253 vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__inv_2
XANTENNA__3968__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3749_ net278 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2012__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2644__A3 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3357__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4632__400 vssd1 vssd1 vccd1 vccd1 _4632__400/HI net400 sky130_fd_sc_hd__conb_1
XANTENNA__2317__C1 team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4123__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2080_ team_10_WB.instance_to_wrap.dispFSM.guesses\[32\] net114 net140 net681 vssd1
+ vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3321__X _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2979__A1_N _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3045__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2982_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] _0837_ net165 vssd1 vssd1 vccd1
+ vccd1 _1489_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_32_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1933_ _0850_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__and2_1
XANTENNA__2812__S net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4652_ net420 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
Xinput30 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
X_1864_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1 vccd1 vccd1
+ _0789_ sky130_fd_sc_hd__inv_2
X_3603_ net277 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4583_ net450 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
Xinput41 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_99_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3534_ net237 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__inv_2
X_3465_ team_10_WB.instance_to_wrap.host_row1\[62\] team_10_WB.instance_to_wrap.dispFSM.msg\[6\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload28_A clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2416_ _1177_ net231 _0849_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__and3b_2
X_3396_ team_10_WB.instance_to_wrap.host_row1\[43\] _1693_ _1770_ _1771_ _1772_ vssd1
+ vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_149_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2347_ _1117_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nand2_1
X_2278_ _0950_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__nor2_1
X_4017_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[1\]
+ net243 vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3036__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4146__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4011__Q team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4296__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input19_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4549__360 vssd1 vssd1 vccd1 vccd1 _4549__360/HI net360 sky130_fd_sc_hd__conb_1
XFILLER_0_155_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2250__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3250_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\] _1608_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__a21o_1
X_3181_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__or4b_1
X_2201_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] _0989_ _0973_ vssd1
+ vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2132_ net214 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0931_ sky130_fd_sc_hd__mux2_1
X_2063_ team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] net109 net135 net678 vssd1
+ vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4019__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1947__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4169__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2965_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\] net161 _1483_ net213
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[12\]
+ sky130_fd_sc_hd__o22a_1
X_4678__433 vssd1 vssd1 vccd1 vccd1 _4678__433/HI net433 sky130_fd_sc_hd__conb_1
X_2896_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\] net153 net121 net616
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[1\]
+ sky130_fd_sc_hd__o22a_1
X_1916_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\] vssd1 vssd1 vccd1 vccd1
+ _0839_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4635_ net403 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4566_ net441 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_25_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3517_ net233 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1953__Y _0875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4497_ net308 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3448_ team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] net170 net169 team_10_WB.instance_to_wrap.dispFSM.msg\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__a22o_1
X_3379_ team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] net173 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[2\]
+ _1756_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__a221o_1
XFILLER_0_169_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1991__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4311__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2750_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ team_10_WB.instance_to_wrap.clock_div.count\[18\] _1365_ vssd1 vssd1 vccd1 vccd1
+ _1372_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_14_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4461__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2681_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4420_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[17\]
+ _0403_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_151_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4351_ clknet_leaf_22_wb_clk_i _0741_ _0340_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[74\]
+ sky130_fd_sc_hd__dfstp_1
X_3302_ _1681_ _1682_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__nand2_1
X_4282_ clknet_leaf_19_wb_clk_i net531 _0271_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3233_ net172 _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3164_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] _1278_ _1568_ _0903_ vssd1 vssd1
+ vccd1 vccd1 _1592_ sky130_fd_sc_hd__a211o_1
X_3095_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] net198 vssd1 vssd1 vccd1
+ vccd1 _1542_ sky130_fd_sc_hd__and2_1
X_2115_ _0916_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_65_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ team_10_WB.instance_to_wrap.dispFSM.guesses\[66\] net111 net137 net693 vssd1
+ vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_105_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3997_ clknet_leaf_27_wb_clk_i _0487_ _0065_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_2948_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] net163 _1478_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[0\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4618_ net389 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_161_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3892__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2879_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net223 vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout111_X net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4549_ net360 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3478__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4334__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4484__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload19 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_23_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3307__A team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3469__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3920_ net268 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3851_ net249 vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2802_ _1409_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__inv_2
X_3782_ net292 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2733_ team_10_WB.instance_to_wrap.clock_div.count\[12\] _1360_ vssd1 vssd1 vccd1
+ vccd1 _1361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2664_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1321_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4207__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4403_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[0\]
+ _0386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2595_ _0908_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__or2_1
X_4334_ clknet_leaf_17_wb_clk_i _0724_ _0323_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[57\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_157_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout206 net208 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_4
Xfanout217 team_10_WB.instance_to_wrap.gamelogic.state\[1\] vssd1 vssd1 vccd1 vccd1
+ net217 sky130_fd_sc_hd__buf_2
Xfanout228 _0846_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
XANTENNA__4357__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4265_ clknet_leaf_5_wb_clk_i _0655_ _0254_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkload10_A clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3216_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] _1626_ vssd1 vssd1 vccd1
+ vccd1 _1628_ sky130_fd_sc_hd__and2_1
X_4196_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[58\]
+ _0185_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[58\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2132__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout273_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3147_ _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__nor2_1
X_3078_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] _1533_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[75\] sky130_fd_sc_hd__mux2_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2029_ net195 _0909_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold260 team_10_WB.instance_to_wrap.dispFSM.guesses\[11\] vssd1 vssd1 vccd1 vccd1
+ net716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_10_WB.instance_to_wrap.clock_div.count\[25\] vssd1 vssd1 vccd1 vccd1
+ net727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\] vssd1 vssd1 vccd1 vccd1
+ net738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2966__A team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2206__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2380_ _0871_ _1088_ _1152_ _1075_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__a32o_1
XANTENNA__3324__X _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4050_ clknet_leaf_14_wb_clk_i _0535_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3001_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\] net164 _1497_ net215
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[34\]
+ sky130_fd_sc_hd__o22a_1
Xinput6 gpio_in[37] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_188_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3903_ net296 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3834_ net272 vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2116__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1955__A team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3765_ net262 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__inv_2
XANTENNA__3393__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2716_ _1171_ _1349_ _1350_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3696_ net246 vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout119_A _0875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2647_ _1307_ _1308_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2578_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] _0898_ _0901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__o2bb2a_1
X_4317_ clknet_leaf_14_wb_clk_i _0707_ _0306_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[40\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3381__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4248_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[4\]
+ _0237_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4179_ clknet_leaf_12_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[41\]
+ _0168_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[41\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_182_Right_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4014__Q team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3384__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4052__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1880_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1 vccd1
+ _0805_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3319__X _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3375__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3550_ net263 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2501_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3481_ team_10_WB.instance_to_wrap.host_row2\[71\] team_10_WB.instance_to_wrap.dispFSM.guesses\[47\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__mux2_1
X_2432_ net194 _1186_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2363_ net228 _0847_ _0853_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__and3b_1
XFILLER_0_138_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4102_ clknet_leaf_24_wb_clk_i _0573_ _0101_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4033_ clknet_leaf_11_wb_clk_i _0518_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2294_ _0859_ _0865_ _1071_ _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout236_A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3817_ net270 vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3748_ net292 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__inv_2
XANTENNA__3366__A2 _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3679_ net272 vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__inv_2
X_4510__321 vssd1 vssd1 vccd1 vccd1 _4510__321/HI net321 sky130_fd_sc_hd__conb_1
XFILLER_0_186_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4075__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4009__Q team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3357__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3315__A team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4418__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2981_ net211 _1485_ _1488_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[23\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1932_ team_10_WB.instance_to_wrap.host_col\[3\] net224 team_10_WB.instance_to_wrap.host_col\[1\]
+ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__or4_2
XFILLER_0_126_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4651_ net419 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
X_1863_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1
+ _0788_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_3602_ net281 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4582_ net449 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
Xinput42 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_99_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3533_ net241 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__inv_2
X_3464_ _1828_ _1831_ _1837_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__o21a_1
X_2415_ net231 _1171_ net458 vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a21oi_1
X_3395_ team_10_WB.instance_to_wrap.host_row1\[51\] _1699_ net179 team_10_WB.instance_to_wrap.host_row2\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4098__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2346_ _0829_ _1121_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _1122_ sky130_fd_sc_hd__a21o_1
X_2277_ _1054_ _1055_ _1058_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__and3b_1
Xclkbuf_2_2__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4016_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[0\]
+ net256 vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4206__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4655__423 vssd1 vssd1 vccd1 vccd1 _4655__423/HI net423 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_167_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2200_ _0919_ _0971_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__a21oi_1
X_3180_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__or4b_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2131_ net134 _0930_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__and2_1
XANTENNA__4390__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2062_ team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] net111 net136 net689 vssd1
+ vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__o22a_1
XFILLER_0_158_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2964_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] net161 _1483_ net214
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[11\]
+ sky130_fd_sc_hd__o22a_1
X_1915_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] vssd1 vssd1 vccd1 vccd1
+ _0838_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2895_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\] net154 net122 net589
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[0\]
+ sky130_fd_sc_hd__o22a_1
X_4634_ net402 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
X_4639__407 vssd1 vssd1 vccd1 vccd1 _4639__407/HI net407 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_155_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4565_ net440 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3516_ net233 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__inv_2
X_4496_ net307 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3447_ team_10_WB.instance_to_wrap.dispFSM.guesses\[21\] net174 net167 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\]
+ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__a22o_1
XANTENNA__2701__A0 team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3378_ team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] _1715_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[66\]
+ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2329_ _0819_ _0849_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] vssd1
+ vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_68_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2018__B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4113__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1991__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1873__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input31_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2471__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2680_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ _1327_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ clknet_leaf_18_wb_clk_i _0740_ _0339_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[73\]
+ sky130_fd_sc_hd__dfstp_1
X_3301_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net210 vssd1 vssd1 vccd1
+ vccd1 _1682_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ clknet_leaf_16_wb_clk_i _0671_ _0270_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_3232_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] _1637_ vssd1 vssd1 vccd1
+ vccd1 _1638_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3163_ _1586_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__xor2_1
X_2114_ team_10_WB.instance_to_wrap.gamelogic.state\[0\] net217 vssd1 vssd1 vccd1
+ vccd1 _0917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3094_ net207 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] net191 _1541_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[83\] sky130_fd_sc_hd__a31o_1
XFILLER_0_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2045_ team_10_WB.instance_to_wrap.dispFSM.guesses\[67\] net110 net138 net640 vssd1
+ vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__o22a_1
XANTENNA__4136__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3996_ clknet_leaf_27_wb_clk_i _0486_ _0064_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2947_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] net163 _1475_ _1476_ _1477_
+ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__o2111ai_4
XANTENNA__4286__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4617_ net388 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2878_ net193 _1462_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[2\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__1973__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4548_ net359 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XANTENNA__2922__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4479_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[36\]
+ _0462_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_5_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2438__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2453__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1868__A team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1964__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1964__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4009__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2211__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3323__A team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4159__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ net272 vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2801_ net230 _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3781_ net263 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_193_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2732_ _1359_ _1360_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[11\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2663_ net513 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\] _1320_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_152_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2594_ _0890_ net226 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\] vssd1
+ vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__a21o_1
X_4402_ clknet_leaf_2_wb_clk_i _0787_ _0385_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\]
+ sky130_fd_sc_hd__dfrtp_4
X_4333_ clknet_leaf_14_wb_clk_i _0723_ _0322_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[56\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_157_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout229 _0018_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_4
X_4571__446 vssd1 vssd1 vccd1 vccd1 net446 _4571__446/LO sky130_fd_sc_hd__conb_1
Xfanout207 team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 net207
+ sky130_fd_sc_hd__clkbuf_4
X_4264_ clknet_leaf_1_wb_clk_i _0654_ _0253_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2380__B2 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout218 team_10_WB.instance_to_wrap.gamelogic.state\[0\] vssd1 vssd1 vccd1 vccd1
+ net218 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3215_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\] _1624_ _1627_ _1611_
+ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4195_ clknet_leaf_12_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[57\]
+ _0184_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[57\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3146_ _1573_ _1574_ _1569_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__a21oi_1
X_3077_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2028_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout266_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3979_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[16\]
+ _0047_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold261 team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] vssd1 vssd1 vccd1 vccd1
+ net717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold250 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\] vssd1 vssd1 vccd1
+ vccd1 net706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold272 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net728 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4301__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2371__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold283 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\] vssd1 vssd1 vccd1 vccd1
+ net739 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3320__B1 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4451__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3387__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3000_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\] net166 _1497_ net216
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[33\]
+ sky130_fd_sc_hd__o22a_1
Xinput7 wb_rst_i vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3902_ net286 vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3833_ net286 vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__inv_2
XANTENNA__3378__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3764_ net292 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2715_ team_10_WB.instance_to_wrap.clock_div.count\[4\] _1347_ team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__a21oi_1
X_3695_ net245 vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2646_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] _0827_ team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__or3_1
XANTENNA__4324__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2577_ _1254_ _1255_ _1260_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4474__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4316_ clknet_leaf_22_wb_clk_i _0706_ _0305_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_4247_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[3\]
+ _0236_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4178_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[40\]
+ _0167_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[40\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout171_X net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3129_ _1557_ _1559_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3369__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3991__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4347__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2500_ net219 net221 net222 net220 vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__or4b_2
X_3480_ team_10_WB.instance_to_wrap.host_row2\[55\] net170 _1848_ _1852_ vssd1 vssd1
+ vccd1 vccd1 _1853_ sky130_fd_sc_hd__a211o_1
X_2431_ net194 _1186_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_94_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2362_ _1091_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__and2b_1
X_4101_ clknet_leaf_24_wb_clk_i _0572_ _0100_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2293_ _0843_ _0846_ net196 _0858_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__nand4b_1
X_4032_ clknet_leaf_13_wb_clk_i _0517_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_1__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2127__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_A _1183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3816_ net252 vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3747_ net260 vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__inv_2
X_3678_ net271 vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2629_ _0807_ _0808_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.blue sky130_fd_sc_hd__nor2_1
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1876__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload7_A clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2980_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] net161 _1488_ net212
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[22\]
+ sky130_fd_sc_hd__o22a_1
X_1931_ net228 _0848_ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1
+ vccd1 _0854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4650_ net418 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_126_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput21 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3601_ net277 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput32 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_we_i vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
X_4581_ net201 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3532_ net254 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__inv_2
X_3463_ team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] net179 _1832_ _1836_ vssd1
+ vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__a211o_1
XANTENNA__2308__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2414_ team_10_WB.instance_to_wrap.clock_div.count\[6\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ _1170_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__or4_2
XFILLER_0_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3394_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net209 _1681_ _1686_
+ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__and4_1
X_2345_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _0870_ _1118_ _1120_
+ _0828_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__a32o_1
X_4533__344 vssd1 vssd1 vccd1 vccd1 _4533__344/HI net344 sky130_fd_sc_hd__conb_1
XFILLER_0_165_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2276_ _0791_ net211 _1050_ _1053_ _1057_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4015_ clknet_leaf_21_wb_clk_i _0503_ net263 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout179_A _1727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2492__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4042__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4192__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2483__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Left_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2214__B net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4517__328 vssd1 vssd1 vccd1 vccd1 _4517__328/HI net328 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_168_Left_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2130_ net213 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0930_ sky130_fd_sc_hd__mux2_1
X_2061_ team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] net110 net138 net679 vssd1
+ vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__o22a_1
XFILLER_0_158_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_177_Left_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3423__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2963_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] net165 _1483_ net215
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[10\]
+ sky130_fd_sc_hd__o22a_1
X_1914_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\] vssd1 vssd1 vccd1 vccd1
+ _0837_ sky130_fd_sc_hd__inv_2
X_4604__378 vssd1 vssd1 vccd1 vccd1 _4604__378/HI net378 sky130_fd_sc_hd__conb_1
X_2894_ net160 net152 vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ net401 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_155_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4564_ net439 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3515_ net233 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__inv_2
XANTENNA__4065__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4495_ net306 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_186_Left_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3446_ team_10_WB.instance_to_wrap.dispFSM.guesses\[77\] _1715_ _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[13\]
+ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3377_ team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] net180 net179 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\]
+ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2328_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\] _0858_ vssd1 vssd1
+ vccd1 vccd1 _1104_ sky130_fd_sc_hd__xor2_1
XANTENNA__2701__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2259_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0798_ _1036_ _1037_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_68_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1976__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4408__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_177_Right_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1991__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2940__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4088__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3327__Y _1707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3300_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _0817_ vssd1 vssd1 vccd1
+ vccd1 _1681_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_187_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ clknet_leaf_16_wb_clk_i _0670_ _0269_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_3231_ _1637_ _1611_ _1636_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and3b_1
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3162_ _0812_ net4 _0906_ _1582_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__and4_1
X_2113_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__nand2b_1
X_3093_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net198 vssd1 vssd1 vccd1
+ vccd1 _1541_ sky130_fd_sc_hd__and2_1
X_2044_ team_10_WB.instance_to_wrap.dispFSM.guesses\[68\] net110 net138 net666 vssd1
+ vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__o22a_1
XFILLER_0_162_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3995_ clknet_leaf_27_wb_clk_i _0485_ _0063_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2946_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\]
+ net163 vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__a41o_1
XANTENNA__3411__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2135__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2877_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] _1461_ vssd1 vssd1 vccd1
+ vccd1 _1462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout211_A team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4616_ net387 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4547_ net358 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
X_4539__350 vssd1 vssd1 vccd1 vccd1 _4539__350/HI net350 sky130_fd_sc_hd__conb_1
XFILLER_0_142_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4478_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[35\]
+ _0461_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\]
+ sky130_fd_sc_hd__dfstp_1
X_3429_ net303 team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _0815_ net209 vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_5_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3478__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2989__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1964__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4380__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3948__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3469__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2429__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3780_ net293 vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__inv_2
X_2800_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[4\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2731_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ _1356_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4401_ clknet_leaf_7_wb_clk_i _0786_ _0384_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_10_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2662_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ _1318_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_152_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2593_ _0910_ _1276_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__nand2_2
X_4332_ clknet_leaf_21_wb_clk_i _0722_ _0321_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout208 team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 net208
+ sky130_fd_sc_hd__clkbuf_2
Xfanout219 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\] vssd1 vssd1 vccd1
+ vccd1 net219 sky130_fd_sc_hd__buf_2
X_4263_ clknet_leaf_1_wb_clk_i _0653_ _0252_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3214_ _1626_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__inv_2
X_4194_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[56\]
+ _0183_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[56\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3145_ _1569_ _1573_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__and3_1
X_3076_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] _1532_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[74\] sky130_fd_sc_hd__mux2_1
XANTENNA__4253__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2027_ _0888_ _0908_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout161_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3978_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[15\]
+ _0046_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2929_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] net151 net120 net682
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[34\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold251 team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] vssd1 vssd1 vccd1 vccd1
+ net707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] vssd1 vssd1 vccd1 vccd1
+ net696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 team_10_WB.instance_to_wrap.clock_div.count\[2\] vssd1 vssd1 vccd1 vccd1
+ net718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\] vssd1 vssd1 vccd1 vccd1
+ net729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\] vssd1 vssd1 vccd1
+ vccd1 net740 sky130_fd_sc_hd__dlygate4sd3_1
X_4617__388 vssd1 vssd1 vccd1 vccd1 _4617__388/HI net388 sky130_fd_sc_hd__conb_1
XANTENNA__3320__B2 team_10_WB.instance_to_wrap.host_row1\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3084__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1879__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4126__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3334__A _1707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
Xclkbuf_2_0__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3340__Y _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3901_ net249 vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3832_ net267 vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3763_ net259 vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2714_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ _1347_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3694_ net245 vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2645_ net1 net158 team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1
+ vccd1 vccd1 _1307_ sky130_fd_sc_hd__and3b_1
XFILLER_0_168_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4401__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4315_ clknet_leaf_15_wb_clk_i _0705_ _0304_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[38\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2576_ net220 net226 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] vssd1
+ vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_113_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4246_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[2\]
+ _0235_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4177_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[2\]
+ _0166_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3128_ _1286_ _1288_ _1291_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__or4b_1
XFILLER_0_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3059_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3066__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4149__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4299__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_140_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2430_ _0993_ _1185_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__and2_2
XANTENNA__3335__Y _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2361_ _1096_ _1131_ _1135_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__and3_1
X_4100_ clknet_leaf_12_wb_clk_i _0571_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_2292_ _0842_ _0866_ _1070_ _0865_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4031_ clknet_leaf_14_wb_clk_i _0516_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2271__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3815_ net253 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
X_3746_ net283 vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__inv_2
XANTENNA__4441__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3677_ net269 vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
XANTENNA__2430__X _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2797__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2628_ _0009_ _0010_ _0008_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2559_ net218 _0952_ _1024_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4229_ clknet_leaf_1_wb_clk_i _0645_ _0218_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3039__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2014__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_X clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4314__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1930_ net225 _0851_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4464__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput11 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_1
XFILLER_0_181_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput22 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3600_ net270 vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__inv_2
X_4580_ net199 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3531_ net254 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3462_ team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] net171 _1833_ _1835_ vssd1
+ vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__a211o_1
X_3393_ team_10_WB.instance_to_wrap.host_row2\[83\] _1701_ net168 team_10_WB.instance_to_wrap.host_row2\[75\]
+ _1769_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__a221o_1
X_2413_ _1167_ _1173_ _1174_ _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__or4_1
X_2344_ _0823_ _1857_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] vssd1 vssd1
+ vccd1 vccd1 _1120_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2275_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] _1056_ vssd1 vssd1
+ vccd1 vccd1 _1057_ sky130_fd_sc_hd__nor2_1
X_4014_ clknet_leaf_21_wb_clk_i _0502_ net258 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[6\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2244__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3729_ net246 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__inv_2
XANTENNA__3981__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4337__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4487__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_178_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2235__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1994__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1893__Y _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_4556__367 vssd1 vssd1 vccd1 vccd1 _4556__367/HI net367 sky130_fd_sc_hd__conb_1
XFILLER_0_185_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2060_ team_10_WB.instance_to_wrap.dispFSM.guesses\[52\] net110 net138 net657 vssd1
+ vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__o22a_1
XFILLER_0_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2962_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\] net162 _1483_ net216 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[9\] sky130_fd_sc_hd__o22a_1
XFILLER_0_173_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1913_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\] vssd1 vssd1 vccd1 vccd1
+ _0836_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4632_ net400 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2893_ net166 net156 vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4500__311 vssd1 vssd1 vccd1 vccd1 _4500__311/HI net311 sky130_fd_sc_hd__conb_1
X_4563_ net374 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
X_4494_ net305 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_155_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3514_ net233 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__inv_2
X_3445_ _0821_ _1819_ _1817_ _1812_ _1807_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkload26_A clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3376_ team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] net174 net170 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\]
+ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout191_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2327_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\] _0854_ vssd1 vssd1
+ vccd1 vccd1 _1103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout289_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2258_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0798_ _0799_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2189_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] net212 vssd1 vssd1 vccd1
+ vccd1 _0978_ sky130_fd_sc_hd__nand2_1
XANTENNA__3398__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3414__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2456__B2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1967__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2392__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ _1633_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__and3_1
X_3161_ team_10_WB.instance_to_wrap.dispFSM.msg\[2\] _0886_ _1274_ _1581_ _1589_ vssd1
+ vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__o32a_1
X_2112_ team_10_WB.instance_to_wrap.dispFSM.guesses\[0\] net114 net141 net645 vssd1
+ vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__o22a_1
X_3092_ net207 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] net191 _1540_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[82\] sky130_fd_sc_hd__a31o_1
X_2043_ net614 net144 net107 net688 vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a22o_1
XANTENNA__3800__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4645__413 vssd1 vssd1 vccd1 vccd1 _4645__413/HI net413 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_105_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3994_ clknet_leaf_27_wb_clk_i _0484_ _0062_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1958__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2945_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] net126 _1474_ vssd1
+ vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2876_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] net223 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_13_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4615_ team_10_WB.instance_to_wrap.gamelogic.red vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
X_4546_ net357 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__4182__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2151__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout204_A team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2922__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4477_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[34\]
+ _0460_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\]
+ sky130_fd_sc_hd__dfstp_1
X_3428_ team_10_WB.instance_to_wrap.host_row1\[53\] net302 _1699_ vssd1 vssd1 vccd1
+ vccd1 _1803_ sky130_fd_sc_hd__o21a_1
XANTENNA_input9_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3332__C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3359_ team_10_WB.instance_to_wrap.host_row1\[41\] _1693_ _1703_ team_10_WB.instance_to_wrap.host_row1\[65\]
+ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout194_X net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_175_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2126__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4055__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2730_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ team_10_WB.instance_to_wrap.clock_div.count\[11\]
+ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_193_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2661_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\] _1319_ vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[0\] sky130_fd_sc_hd__and2b_1
XFILLER_0_81_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4400_ clknet_leaf_2_wb_clk_i _0785_ _0383_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2592_ _0910_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_152_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4331_ clknet_leaf_15_wb_clk_i _0721_ _0320_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[54\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_26_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout209 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\] vssd1 vssd1 vccd1
+ vccd1 net209 sky130_fd_sc_hd__clkbuf_2
X_4262_ clknet_leaf_2_wb_clk_i _0652_ _0251_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_3213_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\] _1621_ vssd1 vssd1 vccd1 vccd1
+ _1626_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4193_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[55\]
+ _0182_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[55\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3144_ _1557_ _1571_ _1572_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__or3_1
X_3075_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2026_ _0888_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3977_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[14\]
+ _0045_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1985__A team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2928_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] net154 net122 net699
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[33\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3396__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _1450_ _1451_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout207_X net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529_ net340 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_170_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold252 team_10_WB.instance_to_wrap.dispFSM.guesses\[70\] vssd1 vssd1 vccd1 vccd1
+ net708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold241 team_10_WB.instance_to_wrap.dispFSM.guesses\[10\] vssd1 vssd1 vccd1 vccd1
+ net697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold230 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\] vssd1 vssd1 vccd1
+ vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] vssd1 vssd1 vccd1
+ vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1 vccd1 vccd1
+ net719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 team_10_WB.instance_to_wrap.dispFSM.guesses\[69\] vssd1 vssd1 vccd1 vccd1
+ net741 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3320__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4078__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3387__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3615__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ net290 vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3831_ net287 vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3762_ net284 vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__inv_2
XANTENNA__3378__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2713_ net655 _1347_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
X_3693_ net246 vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2644_ _0923_ _0947_ _1302_ _0924_ _0922_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[3\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2575_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] net226 net220 vssd1
+ vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4314_ clknet_leaf_21_wb_clk_i net560 _0303_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4220__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4245_ clknet_leaf_32_wb_clk_i net514 _0234_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4176_ clknet_leaf_33_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[1\]
+ _0165_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3127_ _1862_ _1555_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] vssd1
+ vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__a21o_1
XANTENNA__4370__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3058_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _1523_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[65\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2147__Y _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2009_ net219 net220 net221 net222 vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__nor4_2
XTAP_TAPCELL_ROW_120_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3369__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4243__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2360_ _1124_ _1134_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__xor2_1
X_2291_ net5 _0844_ net196 vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__and3_1
XANTENNA__4393__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4030_ clknet_leaf_13_wb_clk_i _0515_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4012__SET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2424__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ net253 vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3745_ net283 vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__inv_2
X_3676_ net291 vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout117_A _0875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2627_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\] _1074_ _1297_ vssd1 vssd1
+ vccd1 vccd1 _0008_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2558_ _1243_ _1247_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nor2_1
X_2489_ net490 _1184_ _1189_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] vssd1
+ vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4228_ clknet_leaf_1_wb_clk_i _0644_ _0217_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4159_ clknet_leaf_29_wb_clk_i _0628_ _0148_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4116__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4266__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2014__A2 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2500__C net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2486__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput34 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
XFILLER_0_181_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput23 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3530_ net241 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3461_ team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] net181 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[70\]
+ _1834_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3392_ team_10_WB.instance_to_wrap.host_row1\[75\] _1708_ net180 team_10_WB.instance_to_wrap.host_row2\[59\]
+ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__a22o_1
X_2412_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2_1
X_2343_ _0870_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__nand2_1
X_2274_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0800_ _1051_ _1052_ _1049_
+ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__a221o_1
X_4013_ clknet_leaf_21_wb_clk_i _0501_ net258 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4139__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2492__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4289__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3441__A1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3441__B2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout234_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2238__A1_N team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3944__RESET_B net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1989_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] net147 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__o22a_1
X_3728_ net250 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__inv_2
X_3659_ net291 vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2704__A0 team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2235__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1994__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1994__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3623__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4567__442 vssd1 vssd1 vccd1 vccd1 net442 _4567__442/LO sky130_fd_sc_hd__conb_1
XANTENNA__4431__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2474__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2961_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\] net165 _1483_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[8\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_173_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1912_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\] vssd1 vssd1 vccd1 vccd1
+ _0835_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2892_ net193 _1471_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_71_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4631_ net399 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
X_4562_ net373 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_181_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4493_ net304 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_155_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2421__B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3513_ net233 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3444_ team_10_WB.instance_to_wrap.host_row2\[45\] net174 net169 team_10_WB.instance_to_wrap.host_row1\[61\]
+ _1818_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkload19_A clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2162__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3375_ team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] net167 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_191_Right_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2326_ _1100_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2257_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] team_10_WB.instance_to_wrap.gamelogic.letter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2188_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net215 vssd1 vssd1 vccd1
+ vccd1 _0977_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3414__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout237_X net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1976__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4304__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4454__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3162__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2456__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2208__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4523__334 vssd1 vssd1 vccd1 vccd1 _4523__334/HI net334 sky130_fd_sc_hd__conb_1
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_187_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3341__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3160_ _0903_ _1588_ net195 vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_146_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3091_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] net198 vssd1 vssd1 vccd1
+ vccd1 _1540_ sky130_fd_sc_hd__and2_1
X_2111_ team_10_WB.instance_to_wrap.dispFSM.guesses\[1\] net109 net135 net691 vssd1
+ vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__o22a_1
Xhold1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe vssd1 vssd1 vccd1 vccd1
+ net457 sky130_fd_sc_hd__dlygate4sd3_1
X_2042_ team_10_WB.instance_to_wrap.dispFSM.guesses\[70\] net115 net141 net702 vssd1
+ vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4610__384 vssd1 vssd1 vccd1 vccd1 _4610__384/HI net384 sky130_fd_sc_hd__conb_1
XFILLER_0_162_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2416__B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3971__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3993_ clknet_leaf_27_wb_clk_i _0483_ _0061_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2944_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] _0831_ net164 vssd1 vssd1
+ vccd1 vccd1 _1475_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2875_ net193 _1460_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[1\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__2432__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4327__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4614_ team_10_WB.instance_to_wrap.gamelogic.green vssd1 vssd1 vccd1 vccd1 net73
+ sky130_fd_sc_hd__clkbuf_1
X_4545_ net356 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_142_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_X clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4476_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[33\]
+ _0459_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4477__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_2__f_wb_clk_i_X clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3427_ team_10_WB.instance_to_wrap.host_row2\[61\] team_10_WB.instance_to_wrap.dispFSM.guesses\[37\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__mux2_1
X_3358_ team_10_WB.instance_to_wrap.host_row2\[41\] net174 _1701_ team_10_WB.instance_to_wrap.host_row2\[81\]
+ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2309_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] _1076_ _1077_
+ net166 vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__a31o_1
X_3289_ _1672_ _1673_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__nor2_1
XANTENNA__2438__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4507__318 vssd1 vssd1 vccd1 vccd1 _4507__318/HI net318 sky130_fd_sc_hd__conb_1
XFILLER_0_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3901__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3994__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2660_ _1307_ _1310_ _1313_ _1317_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2591_ _0908_ _1219_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ clknet_leaf_21_wb_clk_i _0720_ _0319_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4261_ clknet_leaf_0_wb_clk_i _0651_ _0250_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.red
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3212_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\] _1622_ _1625_ vssd1 vssd1
+ vccd1 vccd1 _0536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4192_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[54\]
+ _0181_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[54\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3143_ _1557_ _1572_ _1571_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_173_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3074_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] _1531_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[73\] sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2427__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2025_ net3 _0901_ _0907_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__or3_1
XFILLER_0_174_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3976_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[13\]
+ _0044_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout147_A _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2927_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] net155 net123 net661
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[32\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2858_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\] _1448_ net176
+ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__o21ai_1
X_2789_ _1393_ _1395_ _1396_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__nor4_2
Xhold220 team_10_WB.instance_to_wrap.dispFSM.guesses\[72\] vssd1 vssd1 vccd1 vccd1
+ net676 sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ net339 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_170_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold242 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] vssd1 vssd1 vccd1
+ vccd1 net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] vssd1 vssd1 vccd1 vccd1
+ net709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\] vssd1 vssd1 vccd1 vccd1
+ net687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4459_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[16\]
+ _0442_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\]
+ sky130_fd_sc_hd__dfstp_1
Xhold264 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\] vssd1 vssd1 vccd1
+ vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\] vssd1 vssd1 vccd1 vccd1
+ net742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 team_10_WB.instance_to_wrap.host_row1\[59\] vssd1 vssd1 vccd1 vccd1 net731
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_0_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4172__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529__340 vssd1 vssd1 vccd1 vccd1 _4529__340/HI net340 sky130_fd_sc_hd__conb_1
XFILLER_0_86_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3830_ net271 vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3761_ net283 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2712_ _1347_ _1348_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3692_ net257 vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2643_ _0953_ _1306_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2574_ net221 net226 vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nand2_1
X_4313_ clknet_leaf_18_wb_clk_i _0703_ _0302_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4244_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[0\]
+ _0233_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4175_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[0\]
+ _0164_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3126_ _1286_ _1554_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__nor3_1
XFILLER_0_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3057_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout264_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2008_ net221 _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_120_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3959_ clknet_leaf_31_wb_clk_i _0010_ _0027_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_172_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4045__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4195__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4630__398 vssd1 vssd1 vccd1 vccd1 _4630__398/HI net398 sky130_fd_sc_hd__conb_1
XFILLER_0_185_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2290_ _0842_ _1067_ _0859_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_63_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3813_ net262 vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_72_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2424__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3744_ net264 vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__inv_2
XANTENNA__4068__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3675_ net286 vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2626_ _0828_ _1117_ _1132_ _1235_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2557_ _1239_ _1241_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_81_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2488_ net550 net132 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\] vssd1
+ vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__a22o_1
X_4227_ clknet_leaf_33_wb_clk_i team_10_WB.instance_to_wrap.host_message_reg.next_state
+ _0216_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.Cstate
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4158_ clknet_leaf_31_wb_clk_i net458 _0147_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ sky130_fd_sc_hd__dfrtp_1
X_4089_ clknet_leaf_12_wb_clk_i _0560_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3109_ team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked _0893_ net227 vssd1 vssd1
+ vccd1 vccd1 _1548_ sky130_fd_sc_hd__and3_4
XFILLER_0_167_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2014__A3 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2486__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2238__B1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4210__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4360__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2260__A team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3460_ team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] net175 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[78\]
+ _0821_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__a221o_1
XANTENNA__2961__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3391_ team_10_WB.instance_to_wrap.host_row2\[51\] net170 _1703_ team_10_WB.instance_to_wrap.host_row1\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__a22o_1
X_2411_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__or4b_1
X_2342_ _0820_ _0864_ _0842_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__a21bo_1
X_2273_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _0798_ _0801_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__o22a_1
X_4012_ clknet_leaf_21_wb_clk_i _0500_ net263 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_165_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2477__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2419__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1988_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_119_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3727_ net250 vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__inv_2
XANTENNA__2952__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3658_ net252 vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2609_ _0886_ _1274_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__nor2_1
X_3589_ net260 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_119_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4233__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3432__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4383__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1994__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout190 net192 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2459__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload5_A clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3423__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ net126 _1482_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__nand2_2
X_2891_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] net1 _1227_ vssd1 vssd1 vccd1
+ vccd1 _1471_ sky130_fd_sc_hd__mux2_1
X_1911_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\] vssd1 vssd1 vccd1 vccd1
+ _0834_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4630_ net398 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_146_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4561_ net372 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4492_ clknet_leaf_6_wb_clk_i _0017_ _0475_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_X clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3512_ net232 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__inv_2
X_3443_ team_10_WB.instance_to_wrap.host_row2\[53\] net170 net167 team_10_WB.instance_to_wrap.host_row2\[77\]
+ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__a22o_1
XANTENNA__4106__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _1747_ _1750_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2325_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1858_ vssd1 vssd1 vccd1 vccd1
+ _1101_ sky130_fd_sc_hd__or4b_1
X_2256_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] net216 vssd1 vssd1 vccd1
+ vccd1 _1038_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout177_A _1399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2187_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net215 vssd1 vssd1 vccd1
+ vccd1 _0976_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3414__A2 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4562__373 vssd1 vssd1 vccd1 vccd1 _4562__373/HI net373 sky130_fd_sc_hd__conb_1
XFILLER_0_155_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1967__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3169__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4129__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3634__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4279__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3090_ net205 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] net189 _1539_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[81\] sky130_fd_sc_hd__a31o_1
Xhold2 team_10_WB.instance_to_wrap.keypadFSMHost.strobe vssd1 vssd1 vccd1 vccd1 net458
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2110_ team_10_WB.instance_to_wrap.dispFSM.guesses\[2\] net111 net137 net697 vssd1
+ vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2041_ net585 net144 net107 net597 vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3992_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[29\]
+ _0060_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_2943_ net707 net160 vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1958__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2874_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] _1459_ vssd1 vssd1 vccd1
+ vccd1 _1460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4613_ team_10_WB.instance_to_wrap.blue vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
X_4544_ net355 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_116_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4475_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[32\]
+ _0458_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkload31_A clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3426_ team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.dispFSM.guesses\[69\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout294_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3357_ team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] net170 net169 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__a221o_1
X_2308_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] _1078_ _1083_
+ _1082_ _1079_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__o32a_1
X_3288_ net629 _1671_ net229 vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__o21ai_1
X_2239_ _0796_ net211 _0799_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _1020_
+ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o221a_1
XFILLER_0_165_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4546__357 vssd1 vssd1 vccd1 vccd1 _4546__357/HI net357 sky130_fd_sc_hd__conb_1
XFILLER_0_192_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4421__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input22_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2590_ net195 _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4260_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[3\]
+ _0249_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_3211_ net172 _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__nor2_1
X_4191_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[53\]
+ _0180_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[53\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3142_ _1286_ _1554_ _1556_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__and3b_1
XFILLER_0_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3073_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2024_ _0904_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3975_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[12\]
+ _0043_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2926_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\] net156 net125 net620
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[31\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__4444__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2857_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\] _1448_ vssd1 vssd1
+ vccd1 vccd1 _1450_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2788_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1397_ vssd1 vssd1 vccd1 vccd1
+ _1398_ sky130_fd_sc_hd__or4bb_1
Xhold210 team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] vssd1 vssd1 vccd1 vccd1
+ net666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4527_ net338 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
Xhold243 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\] vssd1 vssd1 vccd1
+ vccd1 net699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] vssd1 vssd1 vccd1 vccd1
+ net677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold232 team_10_WB.instance_to_wrap.dispFSM.guesses\[69\] vssd1 vssd1 vccd1 vccd1
+ net688 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_170_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold276 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\] vssd1 vssd1 vccd1
+ vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 team_10_WB.instance_to_wrap.dispFSM.guesses\[12\] vssd1 vssd1 vccd1 vccd1
+ net721 sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ clknet_leaf_28_wb_clk_i net595 _0441_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold287 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\] vssd1 vssd1 vccd1
+ vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ team_10_WB.instance_to_wrap.host_row1\[44\] _1693_ net173 team_10_WB.instance_to_wrap.host_row2\[84\]
+ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__a22o_1
X_4389_ clknet_leaf_5_wb_clk_i _0774_ _0372_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3069__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_101_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4635__403 vssd1 vssd1 vccd1 vccd1 _4635__403/HI net403 sky130_fd_sc_hd__conb_1
XFILLER_0_121_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3961__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4317__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2528__A _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4681__434 vssd1 vssd1 vccd1 vccd1 _4681__434/HI net434 sky130_fd_sc_hd__conb_1
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4467__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3760_ net278 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2711_ net684 _1345_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3691_ net263 vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2642_ net218 _0952_ _1306_ _0951_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[1\]
+ sky130_fd_sc_hd__a211o_1
X_2573_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\] _1257_ vssd1 vssd1
+ vccd1 vccd1 _1258_ sky130_fd_sc_hd__xnor2_1
X_4312_ clknet_leaf_16_wb_clk_i _0702_ _0301_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4243_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[7\]
+ _0232_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4174_ clknet_leaf_29_wb_clk_i _0643_ _0163_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3125_ _0824_ _1861_ _1555_ _1291_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__a31o_1
X_3056_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] _1522_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\] sky130_fd_sc_hd__mux2_1
XFILLER_0_93_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2007_ net219 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] vssd1 vssd1
+ vccd1 vccd1 _0890_ sky130_fd_sc_hd__or2_1
XANTENNA__2274__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3471__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_186_Right_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3958_ clknet_leaf_33_wb_clk_i _0009_ _0026_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_2909_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\] net153 net121 net700
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[14\]
+ sky130_fd_sc_hd__o22a_1
X_3889_ net282 vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3984__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3732__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_190_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3453__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3089__A team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3812_ net283 vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3743_ net278 vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3674_ net259 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__inv_2
Xoutput101 net183 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
X_2625_ _0010_ _0007_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[1\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3028__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2556_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] _1243_ _1245_
+ _1242_ _1239_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__o221a_1
X_2487_ net498 net133 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1
+ vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__a22o_1
X_4226_ clknet_leaf_17_wb_clk_i net438 _0215_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[101\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4157_ clknet_leaf_31_wb_clk_i net460 _0146_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3108_ net82 net40 net42 vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__and3b_1
X_4088_ clknet_leaf_12_wb_clk_i _0559_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3039_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__mux2_1
XANTENNA__2247__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout162_X net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3444__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2798__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3995__Q team_10_WB.instance_to_wrap.host_col\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2014__A4 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4012__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4162__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2486__A1 team_10_WB.instance_to_wrap.host_row1\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2806__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2238__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput36 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2260__B _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2410_ team_10_WB.instance_to_wrap.clock_div.count\[2\] team_10_WB.instance_to_wrap.clock_div.count\[4\]
+ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or3_1
X_3390_ _1763_ _1765_ _1766_ net303 vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__o31a_1
XFILLER_0_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2341_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _1112_ _1115_ vssd1 vssd1
+ vccd1 vccd1 _1117_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_149_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2272_ _0792_ net214 _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1
+ vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__a22o_1
XANTENNA__3091__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4011_ clknet_leaf_21_wb_clk_i _0499_ net257 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_165_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3426__A0 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4035__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2435__B _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1987_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net150 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout122_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3726_ net250 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__inv_2
XANTENNA__4185__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3657_ net287 vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2165__A0 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2608_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\] _1275_ _1284_ _1289_
+ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
X_3588_ net260 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2539_ team_10_WB.instance_to_wrap.host_col\[3\] _0852_ _1179_ vssd1 vssd1 vccd1
+ vccd1 _0487_ sky130_fd_sc_hd__mux2_1
X_4590__453 vssd1 vssd1 vccd1 vccd1 net453 _4590__453/LO sky130_fd_sc_hd__conb_1
X_4209_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[71\]
+ _0198_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[71\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1979__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout180 _1709_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_4
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2459__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4058__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3408__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2255__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2890_ _1222_ _1470_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[6\]
+ sky130_fd_sc_hd__and2_1
X_1910_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\] vssd1 vssd1 vccd1 vccd1
+ _0833_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4560_ net371 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3511_ net239 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__inv_2
X_4491_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_state _0474_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.Cstate sky130_fd_sc_hd__dfrtp_4
X_3442_ _1800_ _1813_ _1815_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__or4_1
X_3373_ team_10_WB.instance_to_wrap.host_row1\[66\] _1703_ net180 team_10_WB.instance_to_wrap.host_row2\[58\]
+ _1748_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_114_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_166_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net214 vssd1 vssd1 vccd1
+ vccd1 _1037_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2186_ _0822_ _0952_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_wb_clk_i_X clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4689_ net184 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
X_3709_ net236 vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2138__A0 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4200__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4350__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3341__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge vssd1 vssd1 vccd1 vccd1
+ net459 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ team_10_WB.instance_to_wrap.dispFSM.guesses\[72\] net113 net141 team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3991_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[28\]
+ _0059_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2942_ net211 net156 net125 net631 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[47\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net223 vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__or3b_1
XANTENNA__3097__A team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4612_ net386 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
X_4543_ net354 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_142_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4474_ clknet_leaf_28_wb_clk_i net621 _0457_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4223__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload24_A clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3425_ team_10_WB.instance_to_wrap.host_row1\[45\] net302 _1693_ vssd1 vssd1 vccd1
+ vccd1 _1800_ sky130_fd_sc_hd__o21a_1
XANTENNA__2032__B1_N net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3332__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3356_ team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] net167 _1732_ _1734_ vssd1
+ vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__a211o_1
X_3287_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\] _1671_ vssd1 vssd1 vccd1
+ vccd1 _1672_ sky130_fd_sc_hd__and2_1
X_2307_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout287_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2238_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _0804_ _0800_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4373__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3096__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2169_ team_10_WB.instance_to_wrap.correct\[0\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_Left_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Left_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2062__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4246__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_183_Left_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4396__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3210_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ _1621_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__and3_1
X_4190_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[52\]
+ _0179_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[52\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3141_ _1563_ _1570_ _0905_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_192_Left_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3072_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] _1530_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[72\] sky130_fd_sc_hd__mux2_1
XFILLER_0_173_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2023_ _0893_ _0895_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3974_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[11\]
+ _0042_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2925_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\] net153 net121 net674
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[30\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__2443__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2856_ _1448_ _1449_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2787_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__and4b_1
Xhold200 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] vssd1 vssd1 vccd1
+ vccd1 net656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3002__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold211 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\] vssd1 vssd1 vccd1
+ vccd1 net667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4526_ net337 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
Xhold244 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\] vssd1 vssd1 vccd1
+ vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold222 team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] vssd1 vssd1 vccd1 vccd1
+ net678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] vssd1 vssd1 vccd1 vccd1
+ net689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_170_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4457_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[14\]
+ _0440_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\]
+ sky130_fd_sc_hd__dfstp_1
Xhold255 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1
+ net711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\] vssd1 vssd1 vccd1 vccd1
+ net722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] vssd1 vssd1 vccd1 vccd1
+ net733 sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ team_10_WB.instance_to_wrap.host_row1\[52\] _1699_ net167 team_10_WB.instance_to_wrap.host_row2\[76\]
+ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4388_ clknet_leaf_7_wb_clk_i _0773_ _0371_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_input7_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4513__324 vssd1 vssd1 vccd1 vccd1 _4513__324/HI net324 sky130_fd_sc_hd__conb_1
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3339_ _1687_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout192_X net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4119__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2504__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2809__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2710_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__and4_1
X_3690_ net235 vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__inv_2
X_2641_ _0945_ _1305_ _0936_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__a21o_1
X_2572_ net219 net226 vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
X_4311_ clknet_leaf_17_wb_clk_i _0701_ _0300_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4242_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[6\]
+ _0231_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ clknet_leaf_29_wb_clk_i _0642_ _0162_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_3124_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3055_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__mux2_1
XANTENNA__2259__C1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2006_ net219 net220 vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__nor2_1
XANTENNA__2274__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4411__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ clknet_leaf_33_wb_clk_i _0008_ _0025_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2908_ net575 net156 net125 net600 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[13\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3888_ net274 vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4658__426 vssd1 vssd1 vccd1 vccd1 _4658__426/HI net426 sky130_fd_sc_hd__conb_1
X_2839_ _0518_ _1439_ _1436_ _1411_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_115_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4509_ net320 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_131_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4091__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2635__Y _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4434__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3089__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3811_ net262 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4262__Q team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3742_ net292 vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ net287 vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__inv_2
XFILLER_0_179_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2624_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] _1074_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2192__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2192__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2555_ _1246_ _1239_ _1244_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__and3b_1
X_2486_ team_10_WB.instance_to_wrap.host_row1\[48\] net131 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__a221o_1
XANTENNA__3044__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4225_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[87\]
+ _0214_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[87\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4156_ clknet_leaf_27_wb_clk_i _0627_ net255 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked
+ sky130_fd_sc_hd__dfrtp_1
X_3107_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1395_ _1547_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.lcd_en sky130_fd_sc_hd__nor3_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ clknet_leaf_12_wb_clk_i _0558_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2247__A2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3038_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] _1513_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[55\] sky130_fd_sc_hd__mux2_1
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2184__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3951__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4172__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2955__B1 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4307__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4519__330 vssd1 vssd1 vccd1 vccd1 _4519__330/HI net330 sky130_fd_sc_hd__conb_1
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4457__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1997__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1997__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3918__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4606__380 vssd1 vssd1 vccd1 vccd1 _4606__380/HI net380 sky130_fd_sc_hd__conb_1
Xinput15 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3371__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2340_ _1112_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__nand2_1
XANTENNA__2269__A team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2271_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] _0803_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ _1048_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_149_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4010_ clknet_leaf_27_wb_clk_i _0498_ net254 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_74_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3974__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1988__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1988__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4583__450 vssd1 vssd1 vccd1 vccd1 net450 _4583__450/LO sky130_fd_sc_hd__conb_1
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1986_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] _0874_ _0882_ net158 vssd1
+ vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3725_ net267 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3039__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout115_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3656_ net255 vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__inv_2
X_2607_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1288_ _1270_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__or4b_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3587_ net260 vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__inv_2
XANTENNA__3362__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2538_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0840_ _1235_ vssd1 vssd1
+ vccd1 vccd1 _0504_ sky130_fd_sc_hd__a21bo_1
X_4208_ clknet_leaf_12_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[70\]
+ _0197_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[70\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2469_ team_10_WB.instance_to_wrap.host_row1\[58\] net130 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\]
+ _1208_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__a221o_1
XANTENNA__4167__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4139_ clknet_leaf_11_wb_clk_i _0610_ _0138_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3353__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout170 _1702_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_4
Xfanout181 _1709_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout192 _0994_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
XANTENNA__3997__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2459__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2919__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3510_ net239 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4490_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[47\]
+ _0473_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3441_ net180 _1802_ _1809_ net173 vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__a22o_1
XANTENNA__3344__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3372_ team_10_WB.instance_to_wrap.host_row2\[50\] net170 net179 team_10_WB.instance_to_wrap.host_row2\[66\]
+ _1749_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_114_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _1097_ _1098_ _0868_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2254_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net214 vssd1 vssd1 vccd1
+ vccd1 _1036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2185_ net134 _0972_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_69_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4152__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1969_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] net150 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\]
+ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2386__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4688_ net183 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
X_3708_ net234 vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__inv_2
X_3639_ net281 vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2196__X _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_21_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3326__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge vssd1 vssd1 vccd1 vccd1
+ net460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4175__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2301__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2266__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3990_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[27\]
+ _0058_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2941_ team_10_WB.instance_to_wrap.gamelogic.letter\[6\] net155 net123 net656 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[46\] sky130_fd_sc_hd__o22a_1
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ net385 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
X_2872_ net193 _1458_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_84_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4270__Q team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4542_ net353 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4473_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[30\]
+ _0456_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_142_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3424_ team_10_WB.instance_to_wrap.host_row1\[77\] net302 _1708_ vssd1 vssd1 vccd1
+ vccd1 _1799_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4619__390 vssd1 vssd1 vccd1 vccd1 _4619__390/HI net390 sky130_fd_sc_hd__conb_1
XFILLER_0_110_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3355_ team_10_WB.instance_to_wrap.dispFSM.guesses\[65\] _1719_ _1733_ net231 vssd1
+ vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkload17_A clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3286_ net296 _1670_ _1671_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__nor3_1
XFILLER_0_29_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2306_ _0841_ _1073_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__or2_2
X_2237_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _0799_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\]
+ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2168_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__or2_1
X_2099_ team_10_WB.instance_to_wrap.dispFSM.guesses\[21\] net144 net107 net577 vssd1
+ vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4626__394 vssd1 vssd1 vccd1 vccd1 _4626__394/HI net394 sky130_fd_sc_hd__conb_1
XFILLER_0_90_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3020__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4048__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4198__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3140_ _0889_ _0894_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__or2_1
XANTENNA__2522__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3071_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2022_ _0892_ _0896_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2038__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3973_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[10\]
+ _0041_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2924_ net586 net156 net125 net608 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[29\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2855_ net694 _1447_ net176 vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4525_ net336 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
X_2786_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1 _1396_
+ sky130_fd_sc_hd__or3_1
Xhold201 team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] vssd1 vssd1 vccd1 vccd1
+ net657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2210__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3047__S net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold212 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] vssd1 vssd1 vccd1
+ vccd1 net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] vssd1 vssd1 vccd1 vccd1
+ net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] vssd1 vssd1 vccd1 vccd1
+ net679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold256 team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] vssd1 vssd1 vccd1 vccd1
+ net712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 team_10_WB.instance_to_wrap.dispFSM.guesses\[68\] vssd1 vssd1 vccd1 vccd1
+ net701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold278 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] vssd1 vssd1 vccd1
+ vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[13\]
+ _0439_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4340__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold267 team_10_WB.instance_to_wrap.host_row1\[56\] vssd1 vssd1 vccd1 vccd1 net723
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4667__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4387_ clknet_leaf_7_wb_clk_i _0772_ _0370_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ sky130_fd_sc_hd__dfstp_2
X_3407_ net466 net177 _1783_ net229 vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__o211a_1
X_3338_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net210 _1707_ vssd1 vssd1
+ vccd1 vccd1 _1718_ sky130_fd_sc_hd__or3_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4552__363 vssd1 vssd1 vccd1 vccd1 _4552__363/HI net363 sky130_fd_sc_hd__conb_1
XANTENNA__4490__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3269_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\]
+ _1657_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout185_X net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2268__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2825__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_X clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3420__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3480__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4213__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2440__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2991__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2640_ _0926_ net188 vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__nand2_1
XANTENNA__4363__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4495__306 vssd1 vssd1 vccd1 vccd1 _4495__306/HI net306 sky130_fd_sc_hd__conb_1
XFILLER_0_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2571_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] _0898_ vssd1 vssd1
+ vccd1 vccd1 _1256_ sky130_fd_sc_hd__nor2_1
X_4310_ clknet_leaf_19_wb_clk_i _0700_ _0299_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4536__347 vssd1 vssd1 vccd1 vccd1 _4536__347/HI net347 sky130_fd_sc_hd__conb_1
XFILLER_0_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4241_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[5\]
+ _0230_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__1904__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4172_ clknet_leaf_29_wb_clk_i _0641_ _0161_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3123_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] _1288_ _1553_ _0825_
+ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__o31a_1
XFILLER_0_179_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3054_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] _1521_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[63\] sky130_fd_sc_hd__mux2_1
XFILLER_0_179_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ net220 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] net222 vssd1
+ vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__or3_2
XANTENNA__3471__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2454__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3956_ clknet_leaf_33_wb_clk_i _0007_ _0024_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2907_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\] net151 net120 net713
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[12\]
+ sky130_fd_sc_hd__o22a_1
X_3887_ net282 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2838_ _1407_ _0515_ _1426_ _1409_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__o31a_1
X_2769_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[25\]
+ team_10_WB.instance_to_wrap.clock_div.count\[24\] _1380_ vssd1 vssd1 vccd1 vccd1
+ _1384_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4508_ net319 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_131_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4439_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[36\]
+ _0422_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_29_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3462__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4386__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3150__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ net280 vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3741_ net280 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3672_ net259 vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__inv_2
XANTENNA__2964__B2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2623_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1074_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4109__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_112_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2554_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] _1241_ vssd1 vssd1 vccd1
+ vccd1 _1246_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2485_ net525 net130 _1187_ _1215_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4224_ clknet_leaf_12_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[86\]
+ _0213_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[86\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4155_ clknet_leaf_26_wb_clk_i _0626_ _0145_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe
+ sky130_fd_sc_hd__dfrtp_1
X_3106_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ _1546_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] vssd1 vssd1 vccd1 vccd1
+ _1547_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_50_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4086_ clknet_leaf_13_wb_clk_i _0557_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3060__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3037_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__mux2_1
XANTENNA__3444__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4680__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout148_X net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3939_ net255 vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1997__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4363__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput27 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4401__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2269__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2270_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net212 vssd1 vssd1 vccd1
+ vccd1 _1052_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1988__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4273__Q team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1985_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] net146 vssd1 vssd1 vccd1
+ vccd1 _0882_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2937__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3724_ net267 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3655_ net274 vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
XANTENNA__3844__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2606_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] _1287_ vssd1 vssd1
+ vccd1 vccd1 _1288_ sky130_fd_sc_hd__and2_1
X_3586_ net273 vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3055__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2537_ _0871_ _1073_ _1088_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__nand3_1
X_2468_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] net197 vssd1 vssd1
+ vccd1 vccd1 _1208_ sky130_fd_sc_hd__and2_1
XANTENNA__3114__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4207_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[69\]
+ _0196_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[69\] sky130_fd_sc_hd__dfrtp_1
X_2399_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[6\]
+ team_10_WB.instance_to_wrap.clock_div.count\[5\] vssd1 vssd1 vccd1 vccd1 _1162_
+ sky130_fd_sc_hd__or3b_1
X_4138_ clknet_leaf_11_wb_clk_i _0609_ _0137_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3417__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4069_ clknet_leaf_24_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[0\]
+ _0089_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1979__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4226__438 vssd1 vssd1 vccd1 vccd1 net438 _4226__438/LO sky130_fd_sc_hd__conb_1
XANTENNA__4424__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input38_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4358__Q team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout171 _1702_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_4
Xfanout160 _0873_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
Xfanout193 _1222_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XANTENNA__3408__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3041__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3440_ _1707_ _1804_ _1814_ _1717_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3371_ team_10_WB.instance_to_wrap.host_row2\[82\] _1701_ _1708_ team_10_WB.instance_to_wrap.host_row1\[74\]
+ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_114_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _0844_ _0851_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nand2_1
X_2253_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] net213 vssd1 vssd1 vccd1
+ vccd1 _1035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2184_ net134 _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__and2_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4447__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3032__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1968_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] net150 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[27\]
+ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout225_A team_10_WB.instance_to_wrap.host_col\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4687_ net184 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
X_3707_ net234 vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1899_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _0823_ sky130_fd_sc_hd__inv_2
X_3638_ net291 vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__inv_2
X_3569_ net242 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold5 team_10_WB.instance_to_wrap.clock_div.count\[29\] vssd1 vssd1 vccd1 vccd1 net461
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] net156 net125 net686 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[45\] sky130_fd_sc_hd__a22o_1
XFILLER_0_84_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2871_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] _1457_ vssd1 vssd1 vccd1
+ vccd1 _1458_ sky130_fd_sc_hd__mux2_1
X_4610_ net384 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_154_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4541_ net352 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4472_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[29\]
+ _0455_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_3423_ net472 net177 _1798_ net229 vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3354_ team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] net173 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__a22o_1
X_3285_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\]
+ _1666_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2305_ _0841_ _0860_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_1
X_2236_ _0796_ net211 net214 _0797_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__a22o_1
XANTENNA__3096__A3 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2167_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__nand2_1
X_2098_ team_10_WB.instance_to_wrap.dispFSM.guesses\[14\] net115 net141 net709 vssd1
+ vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__o22a_1
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2500__D_N net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3987__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_X clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_98_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_181_Right_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4142__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3070_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _1529_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[71\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4292__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2021_ _0892_ _0894_ net226 vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__or3b_1
XFILLER_0_159_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3972_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[9\]
+ _0040_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2923_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\] net151 net120 net706
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[28\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2854_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ _1444_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__and3_1
X_2785_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\]
+ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4524_ net335 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
Xhold202 team_10_WB.instance_to_wrap.dispFSM.guesses\[20\] vssd1 vssd1 vccd1 vccd1
+ net658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold213 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\] vssd1 vssd1 vccd1
+ vccd1 net669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 team_10_WB.instance_to_wrap.dispFSM.guesses\[43\] vssd1 vssd1 vccd1 vccd1
+ net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 team_10_WB.instance_to_wrap.dispFSM.guesses\[9\] vssd1 vssd1 vccd1 vccd1
+ net691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3852__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold268 team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] vssd1 vssd1 vccd1 vccd1
+ net724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 team_10_WB.instance_to_wrap.dispFSM.guesses\[78\] vssd1 vssd1 vccd1 vccd1
+ net702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\] vssd1 vssd1 vccd1
+ vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[12\]
+ _0438_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_3406_ net231 _1774_ _1782_ _1767_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__a211o_1
Xhold279 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\] vssd1 vssd1 vccd1 vccd1
+ net735 sky130_fd_sc_hd__dlygate4sd3_1
X_4386_ clknet_leaf_2_wb_clk_i _0771_ _0369_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_3337_ _1694_ _1714_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout292_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3063__S net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3268_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ net618 vssd1 vssd1
+ vccd1 vccd1 _1659_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2187__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2219_ net28 net29 vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3199_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] _1392_ vssd1 vssd1 vccd1
+ vccd1 _1617_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3474__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4015__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4165__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2201__A1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input20_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4366__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2268__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2991__A2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2570_ net222 net226 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] vssd1
+ vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4240_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[4\]
+ _0229_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2288__A team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4171_ clknet_leaf_29_wb_clk_i _0640_ _0160_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_184_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3122_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\] _1552_ _0824_ vssd1
+ vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__o21a_1
XANTENNA__4276__Q team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3456__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2259__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3053_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__mux2_1
X_2004_ net299 net3 vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__nand2_1
XANTENNA__4038__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3955_ clknet_leaf_31_wb_clk_i _0006_ _0023_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2906_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\] net153 net121 net647
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[11\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__4188__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3886_ net273 vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout138_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2837_ _1407_ _1436_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2768_ team_10_WB.instance_to_wrap.clock_div.count\[24\] _1382_ net727 vssd1 vssd1
+ vccd1 vccd1 _1383_ sky130_fd_sc_hd__a21oi_1
X_4507_ net318 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_131_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2699_ _0807_ team_10_WB.instance_to_wrap.message_reg.state\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ _1343_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _1344_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4438_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[35\]
+ _0421_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ clknet_leaf_3_wb_clk_i _0754_ _0352_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__3447__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2645__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2110__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4330__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3740_ net292 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4503__314 vssd1 vssd1 vccd1 vccd1 _4503__314/HI net314 sky130_fd_sc_hd__conb_1
XFILLER_0_184_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3671_ net274 vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4480__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2622_ _1116_ _1235_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__nor2_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2553_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_189_Left_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2484_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\] _0991_ vssd1 vssd1 vccd1
+ vccd1 _1215_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4223_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[85\]
+ _0212_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[85\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4154_ clknet_leaf_17_wb_clk_i _0625_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfxtp_1
X_4085_ clknet_leaf_13_wb_clk_i _0556_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3105_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1396_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3036_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _1512_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[54\] sky130_fd_sc_hd__mux2_1
XFILLER_0_179_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2465__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3938_ net271 vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3869_ net260 vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4203__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4353__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput39 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3426__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3371__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4648__416 vssd1 vssd1 vccd1 vccd1 _4648__416/HI net416 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_48_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1984_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] net149 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\]
+ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3723_ net267 vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3654_ net288 vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4226__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2605_ _0888_ _1279_ _0900_ _0899_ _0895_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_70_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3585_ net276 vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3362__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2536_ net515 team_10_WB.instance_to_wrap.buffer.temp_guess\[0\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0505_ sky130_fd_sc_hd__mux2_1
X_2467_ net731 net129 _1207_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__o21a_1
X_4206_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\]
+ _0195_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[68\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4376__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2398_ team_10_WB.instance_to_wrap.clock_div.count\[8\] team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] vssd1 vssd1 vccd1 vccd1 _1161_
+ sky130_fd_sc_hd__or3_1
XANTENNA__3071__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4137_ clknet_leaf_8_wb_clk_i _0608_ _0136_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4068_ clknet_leaf_32_wb_clk_i _0550_ _0088_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_3019_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] net189 vssd1 vssd1 vccd1
+ vccd1 _1504_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3353__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout172 _1612_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
Xfanout150 _0862_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_2
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout194 _0991_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4374__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2919__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4249__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4399__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3344__A2 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ team_10_WB.instance_to_wrap.host_row1\[42\] _1693_ net174 team_10_WB.instance_to_wrap.host_row2\[42\]
+ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _0819_ _0849_ _0851_ _0867_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__or4_1
X_2252_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] _1033_ _1025_ _1027_
+ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_166_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2183_ _0923_ _0947_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4509__320 vssd1 vssd1 vccd1 vccd1 _4509__320/HI net320 sky130_fd_sc_hd__conb_1
XFILLER_0_164_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1967_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] net150 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout120_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3706_ net234 vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4686_ net184 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1898_ net218 vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__inv_2
X_3637_ net269 vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__inv_2
X_3568_ net242 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__inv_2
XANTENNA__4686__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2519_ net503 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] vssd1 vssd1
+ vccd1 vccd1 _0526_ sky130_fd_sc_hd__a22o_1
X_3499_ net238 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3326__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4369__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 team_10_WB.instance_to_wrap.host_row1\[101\] vssd1 vssd1 vccd1 vccd1 net462
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2870_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net223 vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4540_ net351 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_154_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4471_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[28\]
+ _0454_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_3422_ net231 _1788_ _1794_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3353_ team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] net180 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[9\]
+ _1731_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__a221o_1
X_3284_ net728 _1668_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__nor2_1
X_2304_ _0868_ _1080_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__o21a_1
X_2235_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _0800_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__a22o_1
X_2166_ _0936_ _0939_ _0954_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__a21o_1
XANTENNA__4414__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2097_ team_10_WB.instance_to_wrap.dispFSM.guesses\[23\] net145 _0915_ net566 vssd1
+ vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2461__C1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_125_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2999_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\] net163 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[32\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3005__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout123_X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4669_ net431 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_134_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_186_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4094__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4564__439 vssd1 vssd1 vccd1 vccd1 net439 _4564__439/LO sky130_fd_sc_hd__conb_1
XFILLER_0_66_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_X clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_152_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3434__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4437__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2020_ _0899_ _0902_ _0901_ _0896_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3971_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[8\]
+ _0039_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2038__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2922_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\] net155 net123 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[27\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_122_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2853_ _1447_ net176 _1446_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[4\]
+ sky130_fd_sc_hd__and3b_1
X_2784_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4523_ net334 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold214 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\] vssd1 vssd1 vccd1
+ vccd1 net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 team_10_WB.instance_to_wrap.dispFSM.guesses\[40\] vssd1 vssd1 vccd1 vccd1
+ net681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\] vssd1 vssd1 vccd1
+ vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_170_Left_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold247 team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] vssd1 vssd1 vccd1 vccd1
+ net703 sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[11\]
+ _0437_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\]
+ sky130_fd_sc_hd__dfstp_1
Xhold258 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\] vssd1 vssd1 vccd1
+ vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 team_10_WB.instance_to_wrap.clock_div.count\[14\] vssd1 vssd1 vccd1 vccd1
+ net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 team_10_WB.instance_to_wrap.clock_div.count\[8\] vssd1 vssd1 vccd1 vccd1
+ net692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4385_ clknet_leaf_7_wb_clk_i _0770_ _0368_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_clkload22_A clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3405_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\] _1690_ net175 _1775_
+ _1781_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3336_ team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] net167 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[72\]
+ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__a22o_1
XANTENNA__2468__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3267_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ _1658_ vssd1 vssd1
+ vccd1 vccd1 _0561_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout285_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2218_ net25 net24 net27 net26 vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__or4_1
X_3198_ _1393_ _1611_ _1616_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_181_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2149_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] _0943_ vssd1 vssd1 vccd1
+ vccd1 _0944_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3954__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1960__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2268__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3465__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4382__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2569__A net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4170_ clknet_leaf_29_wb_clk_i _0639_ _0159_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_3121_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] _1860_ vssd1 vssd1
+ vccd1 vccd1 _1552_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3052_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] _1520_ net208 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[62\] sky130_fd_sc_hd__mux2_1
XANTENNA__3977__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1920__B net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2003_ team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3954_ clknet_leaf_2_wb_clk_i _0005_ _0022_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_3885_ net277 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__inv_2
X_2905_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\] net151 net120 net720
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[10\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2836_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2195__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2767_ net602 _1382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[24\]
+ sky130_fd_sc_hd__xor2_1
X_4506_ net317 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_131_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3392__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2698_ team_10_WB.instance_to_wrap.message_reg.msg\[0\] team_10_WB.instance_to_wrap.message_reg.msg\[1\]
+ team_10_WB.instance_to_wrap.message_reg.msg\[2\] team_10_WB.instance_to_wrap.message_reg.msg\[3\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4437_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[34\]
+ _0420_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input5_A gpio_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4368_ clknet_leaf_2_wb_clk_i _0753_ _0351_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_4299_ clknet_leaf_15_wb_clk_i _0689_ _0288_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[22\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3319_ _1688_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__and2_4
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4132__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4282__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3773__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2587__A1_N net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4377__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3438__A1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3438__B2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3013__A team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4542__353 vssd1 vssd1 vccd1 vccd1 _4542__353/HI net353 sky130_fd_sc_hd__conb_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3670_ net271 vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2621_ _0006_ _0009_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_112_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2552_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] _1243_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__a21o_1
X_4222_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[84\]
+ _0211_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[84\] sky130_fd_sc_hd__dfrtp_1
X_2483_ net543 net131 _1185_ _1214_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__a22o_1
XANTENNA__4005__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4153_ clknet_leaf_17_wb_clk_i _0624_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4084_ clknet_leaf_13_wb_clk_i _0555_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3104_ team_10_WB.EN_VAL_REG net182 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__or2_1
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3429__A1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3035_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4155__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout150_A _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3937_ net271 vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3868_ net270 vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__inv_2
XANTENNA__4689__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2819_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__or2_1
X_3799_ net279 vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input8_X net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4526__337 vssd1 vssd1 vccd1 vccd1 _4526__337/HI net337 sky130_fd_sc_hd__conb_1
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput29 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_176_Right_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4178__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] _0874_ _0881_ net159 vssd1
+ vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3722_ net267 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3653_ net269 vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2604_ _1268_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\] _1265_ vssd1
+ vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__or3b_2
XFILLER_0_23_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3584_ net253 vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__inv_2
XANTENNA__2570__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2535_ net555 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0506_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2466_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] net198 _1187_
+ _1206_ net130 vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__a221o_1
X_4205_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[67\]
+ _0194_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[67\] sky130_fd_sc_hd__dfrtp_1
X_4136_ clknet_leaf_19_wb_clk_i _0607_ _0135_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_2397_ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ team_10_WB.instance_to_wrap.clock_div.count\[9\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__or4bb_1
XANTENNA__2476__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4067_ clknet_leaf_32_wb_clk_i _0549_ _0087_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3018_ net197 _1503_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[45\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_148_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4320__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 net141 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout173 _1701_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_4
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
Xfanout162 net166 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
Xfanout184 net101 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4470__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 _0885_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_107_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2001__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2320_ _1094_ _1095_ _0869_ _1092_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0798_ _0800_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\]
+ _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2182_ net218 net217 team_10_WB.instance_to_wrap.gamelogic.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _0971_ sky130_fd_sc_hd__or3_1
XFILLER_0_192_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_0_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1966_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0874_ _0878_ net158 vssd1
+ vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3705_ net234 vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__inv_2
X_4685_ net436 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
X_1897_ net299 vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4343__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3636_ net291 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout113_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3567_ net243 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_47_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2518_ _0807_ _0808_ net145 vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__and3_2
X_3498_ net257 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__inv_2
X_2449_ net537 net132 _1191_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4119_ clknet_leaf_9_wb_clk_i _0590_ _0118_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3781__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4385__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4216__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4366__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3014__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4470_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[27\]
+ _0453_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\]
+ sky130_fd_sc_hd__dfstp_1
X_3421_ net179 _1795_ _1796_ net175 _1781_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3352_ team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] net174 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[73\]
+ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__a22o_1
XANTENNA__3691__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2525__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2303_ net224 net225 _0869_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__or3_1
X_3283_ net521 _1666_ _1669_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__o21a_1
X_2234_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] _0805_ vssd1 vssd1 vccd1
+ vccd1 _1016_ sky130_fd_sc_hd__nor2_1
X_2165_ _0942_ _0955_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 _0656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2096_ team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] net114 net141 team_10_WB.instance_to_wrap.dispFSM.guesses\[24\]
+ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_64_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2998_ net126 _1496_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3077__S net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1949_ _0841_ _0871_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_134_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4668_ net182 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout116_X net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3619_ net241 vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__inv_2
X_4599_ net199 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3477__C1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4389__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1963__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3468__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3970_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[7\]
+ _0038_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2921_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\] net151 net120 net648
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[26\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2852_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\]
+ _1442_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__and3_1
X_2783_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4522_ net333 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_31_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold204 team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] vssd1 vssd1 vccd1 vccd1
+ net660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 team_10_WB.instance_to_wrap.dispFSM.guesses\[67\] vssd1 vssd1 vccd1 vccd1
+ net671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\] vssd1 vssd1 vccd1
+ vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[10\]
+ _0436_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3404_ _1777_ _1780_ net177 vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__o21ai_2
Xhold259 team_10_WB.instance_to_wrap.dispFSM.guesses\[19\] vssd1 vssd1 vccd1 vccd1
+ net715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] vssd1 vssd1 vccd1 vccd1
+ net704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] vssd1 vssd1 vccd1 vccd1
+ net693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4384_ clknet_leaf_2_wb_clk_i _0769_ _0367_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_3335_ _1687_ _1714_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__nor2_4
XANTENNA_clkload15_A clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3266_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ net295 vssd1 vssd1
+ vccd1 vccd1 _1658_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2217_ net15 net17 net18 net16 vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__or4bb_1
X_3197_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1616_ sky130_fd_sc_hd__or2_1
XANTENNA__3474__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2148_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nand2_1
XANTENNA__2484__B _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2079_ team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] net109 net135 team_10_WB.instance_to_wrap.dispFSM.guesses\[41\]
+ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__o22a_1
XFILLER_0_165_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_192_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2005__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2198__C1 _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4061__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1960__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2976__B2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4404__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3153__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2288__C team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3120_ net195 _1550_ _1290_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3051_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\]
+ net192 vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__mux2_1
XANTENNA__3456__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2002_ team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3953_ clknet_leaf_23_wb_clk_i _0016_ net243 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2904_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\] net153 net121 net669
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[9\]
+ sky130_fd_sc_hd__o22a_1
X_3884_ net269 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2835_ _1415_ _1426_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2766_ _1381_ _1382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[23\]
+ sky130_fd_sc_hd__nor2_1
X_4505_ net316 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2697_ _1341_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\] vssd1 vssd1
+ vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2b_1
X_4436_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[33\]
+ _0419_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4367_ clknet_leaf_2_wb_clk_i _0752_ _0350_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[4\]
+ sky130_fd_sc_hd__dfstp_2
X_3318_ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4298_ clknet_leaf_20_wb_clk_i _0688_ _0287_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3249_ _1610_ _1647_ net297 vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2495__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3447__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4427__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3383__A1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3383__B2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4393__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2110__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2949__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2620_ _0840_ _0860_ _1295_ _1085_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2551_ _1239_ _1242_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a21boi_1
X_2482_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] net185 vssd1 vssd1 vccd1
+ vccd1 _1214_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_10_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4221_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[83\]
+ _0210_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[83\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3944__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4152_ clknet_leaf_17_wb_clk_i _0623_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfxtp_1
X_4083_ clknet_leaf_13_wb_clk_i _0554_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3429__A2 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3103_ net159 _1302_ net198 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_state
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3034_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _1511_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[53\] sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_179_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3062__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3936_ net268 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout143_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3867_ net276 vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__inv_2
X_2818_ _1410_ _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__nand2_1
X_3798_ net292 vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__inv_2
X_2749_ team_10_WB.instance_to_wrap.clock_div.count\[18\] _1370_ vssd1 vssd1 vccd1
+ vccd1 _1371_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_X clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3117__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
X_4419_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[16\]
+ _0402_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_185_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3053__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1982_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] net146 vssd1 vssd1 vccd1
+ vccd1 _0881_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ net251 vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__inv_2
X_3652_ net294 vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3583_ net276 vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__inv_2
X_2603_ _0016_ _0013_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[1\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2534_ net598 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4122__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2465_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] net194 vssd1 vssd1 vccd1
+ vccd1 _1206_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4204_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[66\]
+ _0193_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[66\] sky130_fd_sc_hd__dfrtp_1
X_2396_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0854_ _1158_ net562 vssd1
+ vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__a22o_1
X_4135_ clknet_leaf_11_wb_clk_i _0606_ _0134_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_4066_ clknet_leaf_32_wb_clk_i _0548_ _0086_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3017_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__mux2_1
XANTENNA__3035__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3919_ net289 vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_189_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout130 _1183_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout174 _1696_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_4
Xfanout141 net142 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout163 net164 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_4
Xfanout152 _1182_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
Xfanout196 _0855_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XFILLER_0_186_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3026__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3019__A team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4145__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4654__422 vssd1 vssd1 vccd1 vccd1 _4654__422/HI net422 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2001__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2001__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _0804_ _1029_ _1031_ vssd1
+ vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4295__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2181_ _0970_ team_10_WB.instance_to_wrap.correct\[0\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3017__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1965_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] net146 vssd1 vssd1 vccd1
+ vccd1 _0878_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3704_ net234 vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2532__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4684_ net183 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1896_ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__inv_2
X_3635_ net288 vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3566_ net243 vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3497_ net256 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__inv_2
X_2517_ team_10_WB.instance_to_wrap.message_reg.state\[1\] net143 _0808_ vssd1 vssd1
+ vccd1 vccd1 _1231_ sky130_fd_sc_hd__o21ai_4
X_2448_ net625 net131 _1187_ _1197_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2379_ _1099_ _1151_ _1135_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_184_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4118_ clknet_leaf_20_wb_clk_i net506 _0117_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_4049_ clknet_leaf_14_wb_clk_i _0534_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4018__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4491__Q team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4168__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4638__406 vssd1 vssd1 vccd1 vccd1 _4638__406/HI net406 sky130_fd_sc_hd__conb_1
XFILLER_0_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input36_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 net70 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3021__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2470__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2470__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1981__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3420_ team_10_WB.instance_to_wrap.host_row2\[44\] team_10_WB.instance_to_wrap.dispFSM.guesses\[20\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3351_ net469 net178 _1730_ net229 vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__o211a_1
X_2302_ _0844_ _0847_ _0853_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o21a_1
X_3282_ net296 _1668_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2233_ _0797_ net214 _0804_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _1014_
+ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o221a_1
X_2164_ _0942_ _0943_ _0957_ _0955_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2095_ team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] net109 net135 net651 vssd1
+ vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_64_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4310__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2461__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2997_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] _1494_ _1495_ vssd1
+ vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3410__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1948_ _0865_ _0870_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nand2b_2
X_4667_ net184 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4460__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1879_ net216 vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3618_ net241 vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__inv_2
X_4598_ net199 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3549_ net257 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__inv_2
XANTENNA__3477__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2945__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3792__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4396__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4333__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload1_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2920_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\] net154 net122 net670
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[25\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_122_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4483__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2851_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] _1444_ vssd1 vssd1
+ vccd1 vccd1 _1446_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_75_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2782_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1392_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4521_ net332 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_142_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4452_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[9\]
+ _0435_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\]
+ sky130_fd_sc_hd__dfstp_1
Xhold205 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\] vssd1 vssd1 vccd1
+ vccd1 net661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\] vssd1 vssd1 vccd1
+ vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3403_ _1685_ _1720_ _1778_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__or4_1
Xhold227 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\] vssd1 vssd1 vccd1 vccd1
+ net683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\] vssd1 vssd1 vccd1
+ vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 team_10_WB.instance_to_wrap.message_reg.state\[0\] vssd1 vssd1 vccd1 vccd1
+ net705 sky130_fd_sc_hd__dlygate4sd3_1
X_4383_ clknet_leaf_4_wb_clk_i _0768_ _0366_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3334_ _1707_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net210 vssd1 vssd1
+ vccd1 vccd1 _1714_ sky130_fd_sc_hd__or3b_2
X_3265_ net295 _1656_ _1657_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__nor3_1
XFILLER_0_147_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3459__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2216_ net21 net20 net23 net22 vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__or4_1
X_3196_ _1391_ _1611_ _1615_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_1_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout173_A _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2147_ _0937_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__nor2_4
X_2078_ team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] net109 net135 net695 vssd1
+ vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__o22a_1
XFILLER_0_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2005__B team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4206__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4570__445 vssd1 vssd1 vccd1 vccd1 net445 _4570__445/LO sky130_fd_sc_hd__conb_1
XANTENNA__4356__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3050_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] _1519_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[61\] sky130_fd_sc_hd__mux2_1
XFILLER_0_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2001_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] net147 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1 vccd1 _0748_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2805__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ clknet_leaf_23_wb_clk_i _0015_ net256 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2903_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\] net155 net123 net673
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[8\]
+ sky130_fd_sc_hd__o22a_1
X_3883_ net276 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__inv_2
X_2834_ _0515_ _1428_ _1435_ _1411_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4504_ net315 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_170_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_17_wb_clk_i_X clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2765_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ _1378_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3392__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2696_ team_10_WB.instance_to_wrap.message_reg.msg\[4\] team_10_WB.instance_to_wrap.message_reg.msg\[5\]
+ team_10_WB.instance_to_wrap.message_reg.msg\[6\] team_10_WB.instance_to_wrap.message_reg.msg\[7\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__mux4_1
X_4435_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[32\]
+ _0418_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_92_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4379__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4366_ clknet_leaf_3_wb_clk_i _0751_ _0349_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3317_ _0815_ net210 _1680_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__or3_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout290_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4297_ clknet_leaf_19_wb_clk_i _0687_ _0286_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_3248_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\] _1608_ vssd1 vssd1 vccd1
+ vccd1 _1647_ sky130_fd_sc_hd__xnor2_1
X_3179_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] _1602_ vssd1 vssd1 vccd1 vccd1
+ _0503_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2016__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3368__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_149_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2550_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__inv_2
X_2481_ team_10_WB.instance_to_wrap.host_row1\[51\] net131 _1187_ _1213_ vssd1 vssd1
+ vccd1 vccd1 _0587_ sky130_fd_sc_hd__a22o_1
X_4220_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[82\]
+ _0209_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[82\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4151_ clknet_leaf_17_wb_clk_i _0622_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_158_Left_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4082_ clknet_leaf_14_wb_clk_i _0553_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3102_ net202 net631 net187 _1545_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[87\]
+ sky130_fd_sc_hd__a31o_1
X_3033_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2535__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4051__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3935_ net291 vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Left_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3866_ net253 vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__inv_2
X_2817_ _0516_ _1409_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nand2_1
X_3797_ net262 vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout303_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2748_ _1369_ _1370_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[17\]
+ sky130_fd_sc_hd__nor2_1
X_2679_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] _1327_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4418_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[15\]
+ _0401_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout301 net6 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_176_Left_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4349_ clknet_leaf_16_wb_clk_i _0739_ _0338_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[72\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2793__X _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_190_Right_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3356__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4074__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1981_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] net148 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_31_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3720_ net251 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3651_ net288 vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3582_ net276 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__inv_2
X_2602_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] _1275_ _1285_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a22o_1
X_2533_ net484 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2464_ team_10_WB.instance_to_wrap.host_row1\[60\] net129 _1194_ _1205_ vssd1 vssd1
+ vccd1 vccd1 _0596_ sky130_fd_sc_hd__o22a_1
X_4203_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[65\]
+ _0192_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[65\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2395_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked net225 _0850_ _1158_ net544
+ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4134_ clknet_leaf_20_wb_clk_i _0605_ _0133_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4417__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4065_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[2\]
+ _0085_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3016_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\] net186 _1502_ net207
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[44\] sky130_fd_sc_hd__o211a_1
XANTENNA_fanout253_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3918_ net289 vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
X_3849_ net272 vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2013__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout131 _1183_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_2
Xfanout120 net124 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_2
X_4532__343 vssd1 vssd1 vccd1 vccd1 _4532__343/HI net343 sky130_fd_sc_hd__conb_1
XANTENNA__4097__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
Xfanout164 net166 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_2
Xfanout142 _0914_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
Xfanout175 _1696_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_2
Xfanout186 _0995_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2001__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4015__RESET_B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2180_ _0936_ _0961_ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1964_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\]
+ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o22a_1
XFILLER_0_141_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4683_ net435 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3703_ net236 vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3634_ net237 vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__inv_2
X_1895_ net225 vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4102__Q team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3565_ net242 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__inv_2
XANTENNA__1953__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2516_ net223 _1225_ _1230_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__a21oi_1
X_3496_ net256 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__inv_2
X_4516__327 vssd1 vssd1 vccd1 vccd1 _4516__327/HI net327 sky130_fd_sc_hd__conb_1
X_2447_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] net194 vssd1 vssd1 vccd1
+ vccd1 _1197_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2378_ _1130_ _1150_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_184_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4117_ clknet_leaf_28_wb_clk_i _0588_ _0116_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_4048_ clknet_leaf_14_wb_clk_i _0533_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4603__377 vssd1 vssd1 vccd1 vccd1 _4603__377/HI net377 sky130_fd_sc_hd__conb_1
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1990__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1990__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_104_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2959__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1863__A team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4012__Q team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold9 net66 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2470__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4112__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1981__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4262__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3350_ _1726_ _1729_ net178 vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__or3b_1
XANTENNA__2930__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2301_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] _1078_ _1076_
+ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__o21a_1
X_3281_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ _1664_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__and3_1
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2232_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net213 vssd1 vssd1 vccd1
+ vccd1 _1014_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2808__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2163_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_88_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2094_ team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] net111 net136 net663 vssd1
+ vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__o22a_1
XFILLER_0_177_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2996_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\] _0838_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ _0839_ net164 vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__a41o_1
XFILLER_0_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1947_ net2 net228 _0858_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nor3_1
X_4666_ net182 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
X_1878_ team_10_WB.instance_to_wrap.gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1
+ _0803_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout216_A team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4597_ net199 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
X_3617_ net237 vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3548_ net263 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3479_ team_10_WB.instance_to_wrap.host_row2\[79\] net167 _1849_ _1851_ vssd1 vssd1
+ vccd1 vccd1 _1852_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_4_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4135__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4285__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2204__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1963__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2979__B1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2850_ _1444_ _1445_ net176 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2781_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_130_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4520_ net331 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_142_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1954__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1954__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\] vssd1 vssd1 vccd1
+ vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[8\]
+ _0434_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold206 team_10_WB.instance_to_wrap.dispFSM.guesses\[73\] vssd1 vssd1 vccd1 vccd1
+ net662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3402_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\] _0815_ net209 _1690_
+ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__a31o_1
Xhold239 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\] vssd1 vssd1 vccd1 vccd1
+ net695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 team_10_WB.instance_to_wrap.clock_div.count\[3\] vssd1 vssd1 vccd1 vccd1
+ net684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4382_ clknet_leaf_7_wb_clk_i _0767_ _0365_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2903__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4008__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3333_ team_10_WB.instance_to_wrap.host_row1\[40\] _1693_ _1700_ _1712_ vssd1 vssd1
+ vccd1 vccd1 _1713_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3264_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\]
+ _1653_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2215_ _0997_ _0998_ _0999_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__or4_1
XFILLER_0_147_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4158__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3195_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\] _1390_ vssd1 vssd1 vccd1
+ vccd1 _1615_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2146_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _0939_ _0940_ vssd1 vssd1
+ vccd1 vccd1 _0941_ sky130_fd_sc_hd__or3_2
XFILLER_0_163_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2077_ team_10_WB.instance_to_wrap.dispFSM.guesses\[35\] net112 net139 net680 vssd1
+ vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2979_ _0800_ _1488_ net158 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[21\]
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_192_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3395__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2005__C net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4649_ net417 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2956__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2370__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4609__383 vssd1 vssd1 vccd1 vccd1 _4609__383/HI net383 sky130_fd_sc_hd__conb_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3386__B1 _1727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4300__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4616__387 vssd1 vssd1 vccd1 vccd1 _4616__387/HI net387 sky130_fd_sc_hd__conb_1
X_2000_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] net147 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 _0749_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__4450__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3951_ clknet_leaf_23_wb_clk_i _0014_ net256 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2902_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\] net157 _1472_ net541
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[7\]
+ sky130_fd_sc_hd__a22o_1
X_3882_ net269 vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2833_ _1423_ _1428_ _0518_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3377__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2764_ team_10_WB.instance_to_wrap.clock_div.count\[23\] _1380_ vssd1 vssd1 vccd1
+ vccd1 _1381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4503_ net314 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_170_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2695_ _1239_ _1246_ _1010_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[2\]
+ sky130_fd_sc_hd__a21bo_1
X_4434_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[31\]
+ _0417_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload20_A clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4365_ clknet_leaf_2_wb_clk_i _0750_ _0348_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[2\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3316_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _1695_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__and3_1
X_4296_ clknet_leaf_16_wb_clk_i _0686_ _0285_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_174_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3247_ _1610_ _1646_ net297 vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a21oi_1
X_3178_ _1277_ _1550_ _1551_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_X clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2129_ net134 _0929_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout169_X net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4323__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4473__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2207__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3359__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2480_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] net194 vssd1 vssd1 vccd1
+ vccd1 _1213_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_130_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4150_ clknet_leaf_17_wb_clk_i _0621_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfxtp_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
X_3101_ _0788_ net202 vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__nor2_1
X_4081_ clknet_leaf_13_wb_clk_i _0552_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3032_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] _1510_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[52\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3990__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3934_ net286 vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__inv_2
X_3865_ net260 vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2816_ _1416_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__or2_1
XANTENNA__4346__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3796_ net292 vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3944__Q team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2747_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ _1365_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__and3_1
X_2678_ net546 _1327_ _1330_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[6\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4417_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[14\]
+ _0400_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout302 net6 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input3_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4348_ clknet_leaf_21_wb_clk_i _0738_ _0337_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4279_ clknet_leaf_22_wb_clk_i _0669_ _0268_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1866__A team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4219__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1980_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] net149 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__o22a_1
XANTENNA__4369__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2246__A1_N team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3650_ net259 vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
X_3581_ net276 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__inv_2
X_2601_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] _1275_ _1285_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2532_ net523 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4202_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\]
+ _0191_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[64\] sky130_fd_sc_hd__dfrtp_1
X_2463_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] net197 team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ net126 vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__a22o_1
X_2394_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _1089_ _1158_ net590 vssd1
+ vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a22o_1
X_4133_ clknet_leaf_3_wb_clk_i _0604_ _0132_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[1\]
+ _0084_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3015_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net191 vssd1 vssd1 vccd1
+ vccd1 _1502_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2491__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629__397 vssd1 vssd1 vccd1 vccd1 _4629__397/HI net397 sky130_fd_sc_hd__conb_1
XANTENNA_fanout246_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3917_ net248 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3848_ net268 vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3779_ net255 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout201_X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_2
Xfanout110 net111 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__buf_2
XANTENNA__2310__A team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_2
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_2
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 net145 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_4
Xfanout176 _1440_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
Xfanout198 _0826_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_166_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1993__C1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4041__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4191__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2473__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3466__A_N team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1963_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _0874_ _0877_ net158 vssd1
+ vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__o211a_1
X_4682_ net183 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
X_3702_ net236 vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__inv_2
X_1894_ team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3633_ net235 vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3564_ net242 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__inv_2
XANTENNA__1953__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3495_ net236 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__inv_2
X_2515_ net223 _1225_ net193 vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__o21ai_1
X_4555__366 vssd1 vssd1 vccd1 vccd1 _4555__366/HI net366 sky130_fd_sc_hd__conb_1
X_2446_ _1187_ _1196_ net572 net129 vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_166_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4116_ clknet_leaf_20_wb_clk_i _0587_ _0115_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2377_ _1126_ _1129_ _1128_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_184_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4047_ clknet_leaf_14_wb_clk_i _0532_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3008__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4064__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2455__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4498__309 vssd1 vssd1 vccd1 vccd1 _4498__309/HI net309 sky130_fd_sc_hd__conb_1
XANTENNA__4407__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1966__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1981__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3280_ _1666_ _1667_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__nor2_1
X_2300_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] _1076_ _1077_
+ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__and3_1
X_2231_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] _0803_ vssd1 vssd1 vccd1
+ vccd1 _1013_ sky130_fd_sc_hd__nor2_1
X_2162_ _0942_ _0944_ _0956_ net704 vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2093_ team_10_WB.instance_to_wrap.dispFSM.guesses\[19\] net113 net139 net677 vssd1
+ vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2995_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ net164 vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__a41o_1
XANTENNA__2125__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4087__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3410__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1946_ _0845_ _0855_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__nand2_1
X_4665_ net430 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_1877_ net214 vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__inv_2
XANTENNA__4113__Q team_10_WB.instance_to_wrap.host_row1\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4596_ net199 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_3616_ net237 vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout111_A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3547_ net257 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__inv_2
X_3478_ team_10_WB.instance_to_wrap.host_row2\[47\] net174 _1708_ team_10_WB.instance_to_wrap.host_row1\[79\]
+ _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2795__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2010__D net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3477__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2429_ net501 net130 net128 net742 vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_145_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__B _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4644__412 vssd1 vssd1 vccd1 vccd1 _4644__412/HI net412 sky130_fd_sc_hd__conb_1
XANTENNA__2437__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2988__B2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_185_Right_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1874__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3165__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3468__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2780_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _1390_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1954__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold207 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\] vssd1 vssd1 vccd1 vccd1
+ net663 sky130_fd_sc_hd__dlygate4sd3_1
X_4450_ clknet_leaf_28_wb_clk_i net542 _0433_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold218 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\] vssd1 vssd1 vccd1
+ vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3401_ net175 net171 net181 vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__or3_1
Xhold229 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] vssd1 vssd1 vccd1
+ vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
X_4381_ clknet_leaf_5_wb_clk_i _0766_ _0364_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3947__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3332_ team_10_WB.instance_to_wrap.host_row1\[72\] _1708_ _1711_ net303 _1706_ vssd1
+ vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3263_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] _1653_ net496 vssd1 vssd1
+ vccd1 vccd1 _1656_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3459__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3194_ _1390_ _1611_ _1614_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and3b_1
X_2214_ net12 net11 net14 net13 vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_1_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ team_10_WB.instance_to_wrap.gamelogic.rights\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__or2_1
X_2076_ team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] net112 net138 net622 vssd1
+ vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout159_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2978_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\] net162 _1488_ net213
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[20\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_192_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3395__A1 team_10_WB.instance_to_wrap.host_row1\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1929_ net225 _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__nor2_1
X_4648_ net416 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_151_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4579_ net200 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4252__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3083__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1875__Y _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3386__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3138__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2212__B net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2897__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] vssd1 vssd1 vccd1
+ vccd1 net546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3950_ clknet_leaf_23_wb_clk_i _0013_ net243 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2901_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\] net153 net121 net623
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[6\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3881_ net277 vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2832_ _1405_ _1433_ _1434_ _1432_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a31o_1
XFILLER_0_170_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2763_ _1379_ _1380_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[22\]
+ sky130_fd_sc_hd__nor2_1
X_4502_ net313 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_170_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2694_ net580 _1009_ _1339_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[1\]
+ sky130_fd_sc_hd__o21bai_1
X_4433_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[30\]
+ _0416_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4125__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4364_ clknet_leaf_3_wb_clk_i _0749_ _0347_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_158_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3315_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ _1682_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__and3_1
X_4295_ clknet_leaf_17_wb_clk_i _0685_ _0284_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2018__C_N net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3246_ _1608_ _1645_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__or2_1
XANTENNA__4275__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3177_ _1283_ _1599_ _1601_ net195 vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2128_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] team_10_WB.instance_to_wrap.buffer.temp_guess\[5\]
+ _0926_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3065__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2059_ net564 net143 net108 net584 vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2040__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3056__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4148__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4298__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
X_3100_ net206 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] net190 _1544_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[86\] sky130_fd_sc_hd__a31o_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
X_4080_ clknet_leaf_13_wb_clk_i _0551_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3031_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__mux2_1
XANTENNA__2893__A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_3_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_34_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3933_ net248 vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3864_ net270 vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2815_ _0514_ _0515_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3795_ net261 vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2746_ team_10_WB.instance_to_wrap.clock_div.count\[17\] _1367_ vssd1 vssd1 vccd1
+ vccd1 _1369_ sky130_fd_sc_hd__nor2_1
XANTENNA__2133__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2677_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] _1327_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4416_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[13\]
+ _0399_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout303 net6 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_4
X_4347_ clknet_leaf_16_wb_clk_i _0737_ _0336_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[70\]
+ sky130_fd_sc_hd__dfstp_1
X_4278_ clknet_leaf_17_wb_clk_i _0668_ _0267_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_3229_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\]
+ _1632_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\] vssd1 vssd1 vccd1 vccd1
+ _1636_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout181_X net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2261__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4440__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1882__A team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3029__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3580_ net270 vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__inv_2
X_2600_ _1270_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2531_ net557 team_10_WB.instance_to_wrap.buffer.temp_guess\[5\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0510_ sky130_fd_sc_hd__mux2_1
X_4201_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[63\]
+ _0190_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[63\] sky130_fd_sc_hd__dfrtp_1
X_2462_ net467 net130 _1204_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a21o_1
X_2393_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _1093_ _1158_ net563 vssd1
+ vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a22o_1
X_4132_ clknet_leaf_10_wb_clk_i _0603_ _0131_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_4063_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[0\]
+ _0083_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_155_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3014_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\] net186 _1501_ net205
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\] sky130_fd_sc_hd__o211a_1
XANTENNA__4313__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3916_ net290 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout141_A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4116__Q team_10_WB.instance_to_wrap.host_row1\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout239_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3847_ net288 vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__inv_2
XANTENNA__4463__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3778_ net281 vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2729_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ _1358_ _1177_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout122 net123 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_2
Xfanout111 net116 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_4
Xfanout133 _1183_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
Xfanout155 _1182_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net145 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout177 _1399_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
Xfanout199 net201 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
Xfanout188 net192 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
Xfanout166 _0872_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1877__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3980__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4336__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_X clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2473__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4661__429 vssd1 vssd1 vccd1 vccd1 _4661__429/HI net429 sky130_fd_sc_hd__conb_1
XFILLER_0_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4486__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1962_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] net146 vssd1 vssd1 vccd1
+ vccd1 _0877_ sky130_fd_sc_hd__or2_1
X_4681_ net434 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1893_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\] vssd1 vssd1 vccd1 vccd1
+ _0817_ sky130_fd_sc_hd__inv_2
X_3701_ net236 vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3632_ net235 vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3563_ net242 vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__inv_2
X_2514_ _1226_ _1229_ net193 vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__and3b_1
X_3494_ net245 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2445_ _0836_ net194 vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4115_ clknet_leaf_10_wb_clk_i _0586_ _0114_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_2376_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] _1084_ _1148_
+ _1149_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout189_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ clknet_leaf_14_wb_clk_i _0531_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4566__441 vssd1 vssd1 vccd1 vccd1 net441 _4566__441/LO sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3413__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4209__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4359__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3404__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3327__A team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2930__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2230_ _0822_ net217 team_10_WB.instance_to_wrap.gamelogic.state\[2\] _0988_ team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__a311o_1
X_2161_ _0942_ _0943_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_88_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4589__452 vssd1 vssd1 vccd1 vccd1 net452 _4589__452/LO sky130_fd_sc_hd__conb_1
X_2092_ team_10_WB.instance_to_wrap.dispFSM.guesses\[20\] net113 net139 net690 vssd1
+ vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__o22a_1
XFILLER_0_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2446__B2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2994_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] net160 vssd1 vssd1 vccd1
+ vccd1 _1493_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1945_ _0845_ net196 vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__and2_1
X_4522__333 vssd1 vssd1 vccd1 vccd1 _4522__333/HI net333 sky130_fd_sc_hd__conb_1
XANTENNA__1957__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4664_ net183 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
X_1876_ net213 vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4595_ net201 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_3615_ net237 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__inv_2
X_3546_ net262 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3477_ team_10_WB.instance_to_wrap.host_row2\[87\] net173 net180 team_10_WB.instance_to_wrap.host_row2\[63\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__a221o_1
XANTENNA__2134__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2428_ net188 _1185_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2359_ _1124_ _1134_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4029_ clknet_leaf_13_wb_clk_i _0514_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_104_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4031__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4181__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input34_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4506__317 vssd1 vssd1 vccd1 vccd1 _4506__317/HI net317 sky130_fd_sc_hd__conb_1
XFILLER_0_127_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold208 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\] vssd1 vssd1 vccd1
+ vccd1 net664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3328__Y _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_44_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4380_ clknet_leaf_7_wb_clk_i _0765_ _0363_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_133_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3400_ _1686_ _1698_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__or3_1
Xhold219 team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] vssd1 vssd1 vccd1 vccd1
+ net675 sky130_fd_sc_hd__dlygate4sd3_1
X_3331_ team_10_WB.instance_to_wrap.host_row2\[56\] net180 net168 team_10_WB.instance_to_wrap.host_row2\[72\]
+ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__a22o_1
XANTENNA__2903__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3262_ net613 _1653_ _1655_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__o21a_1
X_3193_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _1614_
+ sky130_fd_sc_hd__a21o_1
X_2213_ net39 net38 net10 net9 vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__or4_1
X_2144_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2075_ team_10_WB.instance_to_wrap.dispFSM.guesses\[45\] net143 net108 net559 vssd1
+ vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__a22o_1
XANTENNA__4054__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3092__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2977_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] net161 _1488_ net214
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[19\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_192_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3395__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout221_A team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1928_ team_10_WB.instance_to_wrap.host_col\[3\] net224 vssd1 vssd1 vccd1 vccd1 _0851_
+ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_62_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4647_ net415 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_188_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4578_ net200 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_3529_ net254 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_71_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_27_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3386__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold80 team_10_WB.instance_to_wrap.clock_div.count\[0\] vssd1 vssd1 vccd1 vccd1 net536
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4077__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold91 team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] vssd1 vssd1 vccd1 vccd1 net547
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2900_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\] net157 net125 net480
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3880_ net269 vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2831_ _1430_ _1431_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__or2_1
XANTENNA__3377__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2762_ team_10_WB.instance_to_wrap.clock_div.count\[21\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ team_10_WB.instance_to_wrap.clock_div.count\[22\] _1374_ vssd1 vssd1 vccd1 vccd1
+ _1380_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4501_ net312 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4432_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[29\]
+ _0415_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_2693_ _1009_ _1238_ _1339_ _1340_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[0\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4363_ clknet_leaf_3_wb_clk_i _0748_ _0346_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3314_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__nand2_2
X_4294_ clknet_leaf_18_wb_clk_i _0684_ _0283_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_3245_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _1645_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3176_ _1582_ _1600_ _0906_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2127_ net134 _0928_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2058_ team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] net114 net140 net703 vssd1
+ vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2812__A1 _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3368__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3359__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2567__B1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
X_3030_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] _1509_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[51\] sky130_fd_sc_hd__mux2_1
XFILLER_0_144_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3932_ net290 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_34_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3863_ net260 vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__inv_2
X_2814_ _1413_ _1418_ _1416_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3794_ net279 vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2745_ _1367_ _1368_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[16\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4402__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2676_ _1318_ _1328_ _1329_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[5\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_41_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4415_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[12\]
+ _0398_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4346_ clknet_leaf_20_wb_clk_i _0736_ _0335_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[69\]
+ sky130_fd_sc_hd__dfrtp_1
X_4277_ clknet_leaf_16_wb_clk_i _0667_ _0266_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4392__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3228_ net639 _1633_ _1635_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__o21a_1
XANTENNA__2089__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout174_X net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3159_ _1586_ _1587_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_16_wb_clk_i_X clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4115__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2234__A team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4265__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2530_ net470 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0511_ sky130_fd_sc_hd__mux2_1
X_2461_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] net203 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ _1189_ net129 vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__o221a_1
X_4200_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[62\]
+ _0189_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[62\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2392_ net2 net581 _1158_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4131_ clknet_leaf_10_wb_clk_i _0602_ _0130_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_4062_ clknet_leaf_14_wb_clk_i _0547_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3013_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] net189 vssd1 vssd1 vccd1
+ vccd1 _1501_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3915_ net254 vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3440__A1 _1707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3440__B2 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3846_ net286 vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3777_ net284 vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2728_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ vssd1 vssd1 vccd1
+ vccd1 _1358_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout301_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2659_ _1310_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__nand2_2
Xfanout112 net116 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
X_4329_ clknet_leaf_19_wb_clk_i _0719_ _0318_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_2
Xfanout145 _0912_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_2
Xfanout134 _0919_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
Xfanout178 _1399_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
Xfanout167 _1710_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4138__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4288__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3431__A1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2473__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1961_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[32\]
+ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__o22a_1
XANTENNA__3422__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3700_ net235 vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ net184 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
X_1892_ team_10_WB.instance_to_wrap.lcdPlayer.currentState\[0\] vssd1 vssd1 vccd1
+ vccd1 _0816_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1984__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1984__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3631_ net247 vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3347__X _1727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3562_ net242 vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2513_ net223 _1225_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] vssd1
+ vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3493_ net235 vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2444_ net606 net132 _1185_ _1195_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__a22o_1
X_2375_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2161__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4114_ clknet_leaf_20_wb_clk_i _0585_ _0113_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_4045_ clknet_leaf_14_wb_clk_i _0530_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2449__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2139__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2464__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4430__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout251_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3829_ net247 vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2455__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1966__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3327__B _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4303__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4453__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _0936_ _0941_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__a21o_1
X_2091_ net737 net144 net107 net583 vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_183_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2993_ net729 net160 _1492_ net211 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[31\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1944_ _0858_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__or2_1
X_4663_ net183 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
X_4561__372 vssd1 vssd1 vccd1 vccd1 _4561__372/HI net372 sky130_fd_sc_hd__conb_1
XFILLER_0_153_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3614_ net237 vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__inv_2
X_1875_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1 vccd1
+ _0800_ sky130_fd_sc_hd__inv_2
X_4594_ net199 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2422__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3545_ net263 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__inv_2
X_3476_ team_10_WB.instance_to_wrap.host_row1\[55\] _1699_ net169 team_10_WB.instance_to_wrap.host_row1\[63\]
+ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__a22o_1
X_2427_ net185 _1186_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nor2_1
XANTENNA__3331__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2358_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1133_ _1132_ _1117_
+ _1100_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_193_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2289_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4028_ clknet_leaf_13_wb_clk_i _0513_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2437__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3970__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4326__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4476__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input27_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4545__356 vssd1 vssd1 vccd1 vccd1 _4545__356/HI net356 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_26_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3389__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold209 team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] vssd1 vssd1 vccd1 vccd1
+ net665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3330_ _1683_ _1687_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3261_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] _1653_ net295 vssd1 vssd1
+ vccd1 vccd1 _1655_ sky130_fd_sc_hd__a21oi_1
X_3192_ _1389_ _1611_ _1613_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__and3_1
X_2212_ net19 net8 net33 net30 vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__or4_1
XFILLER_0_147_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2143_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.correct\[0\]
+ team_10_WB.instance_to_wrap.correct\[2\] vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2074_ team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] net115 net141 net733 vssd1
+ vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__o22a_1
XANTENNA__3993__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4349__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2976_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\] net161 _1488_ net215
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[18\]
+ sky130_fd_sc_hd__o22a_1
X_1927_ net228 _0848_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout214_A team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4646_ net414 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_188_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4577_ net199 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_151_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3528_ net233 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__inv_2
X_3459_ team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] net173 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__a22o_1
XANTENNA__3430__B _0817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2997__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2897__A2 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold70 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] vssd1 vssd1 vccd1 vccd1
+ net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_10_WB.instance_to_wrap.host_row1\[67\] vssd1 vssd1 vccd1 vccd1 net537
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3621__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 _0512_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2830_ _1430_ _1431_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3339__Y _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2761_ team_10_WB.instance_to_wrap.clock_div.count\[22\] _1378_ vssd1 vssd1 vccd1
+ vccd1 _1379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4500_ net311 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2692_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] _1241_ vssd1 vssd1
+ vccd1 vccd1 _1340_ sky130_fd_sc_hd__or2_1
XANTENNA_1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4431_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[28\]
+ _0414_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4634__402 vssd1 vssd1 vccd1 vccd1 _4634__402/HI net402 sky130_fd_sc_hd__conb_1
X_4362_ clknet_leaf_11_wb_clk_i _0747_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_4293_ clknet_leaf_16_wb_clk_i _0683_ _0282_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_3313_ net210 _1686_ _1688_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__and4b_4
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3244_ _1610_ _1644_ net296 vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3175_ _0887_ _0894_ _0891_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2126_ net212 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout164_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4171__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2057_ net624 net144 net107 net627 vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2959_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] _1480_ _1481_ vssd1
+ vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2576__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629_ net397 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_102_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1896__A team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3616__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4044__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_169_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4194__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3931_ net254 vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3862_ net270 vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__inv_2
X_2813_ _1415_ _1417_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3793_ net279 vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2744_ team_10_WB.instance_to_wrap.clock_div.count\[16\] _1365_ _1177_ vssd1 vssd1
+ vccd1 vccd1 _1368_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2675_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\]
+ _1321_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\] vssd1 vssd1 vccd1
+ vccd1 _1329_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4414_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[11\]
+ _0397_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4345_ clknet_leaf_18_wb_clk_i _0735_ _0334_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4276_ clknet_leaf_33_wb_clk_i _0666_ _0265_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3227_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] _1633_ net172 vssd1
+ vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout281_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2494__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3158_ _1560_ _1585_ _1584_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_178_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2109_ team_10_WB.instance_to_wrap.dispFSM.guesses\[3\] net112 net139 net716 vssd1
+ vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout167_X net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3089_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] net198 vssd1 vssd1 vccd1
+ vccd1 _1539_ sky130_fd_sc_hd__and2_1
XFILLER_0_193_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4067__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2994__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1897__Y _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1996__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2460_ net478 net129 _1203_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4130_ clknet_leaf_19_wb_clk_i _0601_ _0129_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_2391_ net532 _1158_ _1159_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4061_ clknet_leaf_15_wb_clk_i _0546_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3012_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\] net185 _1500_ net204
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[42\] sky130_fd_sc_hd__o211a_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3914_ net272 vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__inv_2
XANTENNA__2425__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3845_ net252 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout127_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3776_ net278 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2727_ _1180_ _1355_ _1357_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[9\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__2951__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_189_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2658_ net193 _1234_ _1225_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__o21bai_2
Xfanout113 net116 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2589_ _1272_ _1273_ _0902_ _0908_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__2703__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4328_ clknet_leaf_17_wb_clk_i _0718_ _0317_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[51\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout124 _1473_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_2
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
Xfanout146 net147 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_148_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout168 _1710_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
Xfanout179 _1727_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_4
XANTENNA_input1_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _1181_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
X_4259_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[2\]
+ _0248_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2942__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_155_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3407__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4232__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_164_Left_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1960_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\]
+ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__o22a_1
XFILLER_0_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1891_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] vssd1 vssd1 vccd1 vccd1
+ _0815_ sky130_fd_sc_hd__inv_2
XANTENNA__4382__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3630_ net248 vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3561_ net242 vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_180_Right_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2512_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] _1226_ _1228_ vssd1
+ vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3492_ net235 vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_173_Left_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2443_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net186 vssd1 vssd1 vccd1
+ vccd1 _1195_ sky130_fd_sc_hd__or2_1
X_2374_ _0871_ _1147_ _1087_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a21oi_1
X_4113_ clknet_leaf_10_wb_clk_i _0584_ _0112_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4044_ clknet_leaf_14_wb_clk_i _0529_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3110__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_182_Left_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3413__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout244_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3828_ net287 vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3759_ net279 vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_191_Left_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4105__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4255__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3624__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2090_ team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] net115 net141 net665 vssd1
+ vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_88_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2527__X _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2992_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net165 _1491_ net212
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[30\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1943_ _0844_ net196 vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__and2_1
X_4662_ net182 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
XANTENNA__1957__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1874_ net212 vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3613_ net241 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4593_ net199 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4128__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3544_ net262 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__inv_2
X_3475_ team_10_WB.instance_to_wrap.host_row1\[47\] _1693_ _1703_ team_10_WB.instance_to_wrap.host_row1\[71\]
+ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkload29_A clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2426_ _0993_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__nor2_2
XANTENNA__3534__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4278__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout194_A _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2357_ _0823_ _0828_ _1859_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2288_ team_10_WB.instance_to_wrap.host_col\[3\] net225 team_10_WB.instance_to_wrap.host_col\[0\]
+ net224 vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__or4b_2
X_4027_ clknet_leaf_33_wb_clk_i net548 _0074_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4651__419 vssd1 vssd1 vccd1 vccd1 _4651__419/HI net419 sky130_fd_sc_hd__conb_1
XFILLER_0_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3086__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4420__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3260_ net463 _1651_ _1654_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__o21a_1
X_3191_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2211_ net35 net34 net37 net36 vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__or4_1
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2142_ _0916_ _0935_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2073_ net568 net143 net108 net628 vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3092__A3 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2975_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\] net161 _1488_ net216
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[17\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1926_ net228 _0848_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__nor2_1
X_4645_ net413 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4576_ net201 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout207_A team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3527_ net232 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__inv_2
X_3458_ team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] net168 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[14\]
+ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__a22o_1
X_3389_ team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] _1701_ net181 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\]
+ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__a22o_1
X_2409_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout197_X net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3068__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4443__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3174__A team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4512__323 vssd1 vssd1 vccd1 vccd1 _4512__323/HI net323 sky130_fd_sc_hd__conb_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold71 team_10_WB.instance_to_wrap.host_row1\[77\] vssd1 vssd1 vccd1 vccd1 net527
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked vssd1 vssd1 vccd1 vccd1
+ net538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 _0505_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold93 team_10_WB.instance_to_wrap.host_row1\[63\] vssd1 vssd1 vccd1 vccd1 net549
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2034__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2760_ _1377_ _1378_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[21\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2691_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] _1246_ _1238_ vssd1
+ vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__a21oi_1
X_4430_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[27\]
+ _0413_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4361_ clknet_leaf_11_wb_clk_i _0004_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3312_ _1691_ _1692_ net283 vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__a21oi_1
X_4292_ clknet_leaf_19_wb_clk_i net567 _0281_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3243_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3960__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3174_ team_10_WB.instance_to_wrap.dispFSM.msg\[6\] _1550_ vssd1 vssd1 vccd1 vccd1
+ _1599_ sky130_fd_sc_hd__or2_1
XANTENNA__3023__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2125_ net134 _0927_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__and2_1
XANTENNA__4316__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2428__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2056_ team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] net115 net140 net654 vssd1
+ vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_37_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2273__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3470__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4466__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2958_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] _0832_ net165 vssd1 vssd1 vccd1
+ vccd1 _1481_ sky130_fd_sc_hd__a41o_1
XFILLER_0_161_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1909_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\] vssd1 vssd1 vccd1 vccd1
+ _0832_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4628_ net396 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2889_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] net1 _1469_ vssd1 vssd1 vccd1
+ vccd1 _1470_ sky130_fd_sc_hd__mux2_1
X_4559_ net370 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3461__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4657__425 vssd1 vssd1 vccd1 vccd1 _4657__425/HI net425 sky130_fd_sc_hd__conb_1
XFILLER_0_152_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2801__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3983__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_169_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4339__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4489__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3930_ net271 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3452__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3861_ net274 vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2812_ _0816_ _0817_ net178 vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3792_ net264 vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2743_ team_10_WB.instance_to_wrap.clock_div.count\[15\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ _1364_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2674_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2430__B _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4413_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[10\]
+ _0396_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_4344_ clknet_leaf_18_wb_clk_i _0734_ _0333_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[67\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_185_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4275_ clknet_leaf_2_wb_clk_i _0665_ _0264_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkload11_A clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3226_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1632_ _1634_ vssd1
+ vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout274_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3157_ _1560_ _1584_ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2108_ team_10_WB.instance_to_wrap.dispFSM.guesses\[4\] net112 net139 net721 vssd1
+ vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__o22a_1
X_3088_ net206 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] net190 _1538_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[80\] sky130_fd_sc_hd__a31o_1
XFILLER_0_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2039_ team_10_WB.instance_to_wrap.dispFSM.guesses\[73\] net111 net136 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_59_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3443__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2237__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2237__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4011__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3627__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4161__CLK clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2390_ _0858_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__nor2_1
X_4060_ clknet_leaf_14_wb_clk_i _0545_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3011_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] net188 vssd1 vssd1 vccd1
+ vccd1 _1500_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3425__B1 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3913_ net288 vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__inv_2
XANTENNA__2425__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3844_ net289 vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__inv_2
XANTENNA__1987__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3775_ net277 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2726_ _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2657_ net193 _1225_ _1227_ _1234_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[2\]
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_189_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2588_ _0898_ _0901_ _0907_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__and3_1
Xfanout114 net115 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_2
Xfanout136 net137 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
X_4327_ clknet_leaf_22_wb_clk_i _0717_ _0316_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[50\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout125 _1472_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
Xfanout147 _0862_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_4
Xfanout169 _1704_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_4
X_4258_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[1\]
+ _0247_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout158 net160 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
X_3209_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] _1621_ _1623_ vssd1 vssd1
+ vccd1 vccd1 _0535_ sky130_fd_sc_hd__o21a_1
X_4189_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[51\]
+ _0178_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[51\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3416__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4184__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\] vssd1 vssd1 vccd1
+ vccd1 net646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3910__A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1969__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1890_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ _0814_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3560_ net242 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2511_ _1225_ _1227_ net193 vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a21boi_1
X_3491_ net237 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2442_ net512 net133 net127 net738 vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3343__C1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2373_ _1137_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__or2_1
X_4112_ clknet_leaf_19_wb_clk_i _0583_ _0111_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4043_ clknet_leaf_14_wb_clk_i _0528_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4057__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3031__S net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout237_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3827_ net247 vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3758_ net293 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2709_ _1345_ _1346_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
X_3689_ net236 vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__inv_2
X_4573__448 vssd1 vssd1 vccd1 vccd1 net448 _4573__448/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_7_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2128__A0 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2256__A team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2991_ net601 net160 _1492_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[29\] sky130_fd_sc_hd__a22o_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1942_ _0819_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__nand2_1
X_4661_ net429 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
X_1873_ net211 vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3612_ net277 vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4592_ net455 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3543_ net263 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__inv_2
X_3474_ team_10_WB.instance_to_wrap.dispFSM.guesses\[31\] net170 net167 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\]
+ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2425_ net197 _0942_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3331__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2356_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1119_ vssd1 vssd1 vccd1
+ vccd1 _1132_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout187_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3550__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2287_ _1064_ _1063_ team_10_WB.instance_to_wrap.gamelogic.rights\[0\] vssd1 vssd1
+ vccd1 vccd1 _0644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4026_ clknet_leaf_0_wb_clk_i net471 _0073_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2070__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4222__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4372__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3389__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3338__C _1707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2210_ _0806_ _0996_ net194 _0945_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__a2bb2o_1
X_3190_ net473 net172 vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2141_ _0916_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nor2_1
X_2072_ team_10_WB.instance_to_wrap.dispFSM.guesses\[40\] net114 net140 net726 vssd1
+ vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2974_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] net161 _1488_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[16\]
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_6_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_1925_ net2 net3 net299 vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__o21ba_1
X_4644_ net412 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_71_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4575_ net200 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3001__B2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4245__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3526_ net232 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__inv_2
XANTENNA__3545__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4395__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3457_ team_10_WB.instance_to_wrap.host_row1\[78\] _1708_ _1829_ _1830_ vssd1 vssd1
+ vccd1 vccd1 _1831_ sky130_fd_sc_hd__a211o_1
X_3388_ team_10_WB.instance_to_wrap.dispFSM.guesses\[75\] _1715_ _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[11\]
+ _1764_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__a221o_1
X_2408_ _1164_ _1167_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__nor3_1
X_2339_ _1110_ _1111_ _1113_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ clknet_leaf_23_wb_clk_i _0497_ net257 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ sky130_fd_sc_hd__dfstp_2
XPHY_EDGE_ROW_40_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4551__362 vssd1 vssd1 vccd1 vccd1 _4551__362/HI net362 sky130_fd_sc_hd__conb_1
XANTENNA_input32_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 _0589_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net71 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] vssd1 vssd1 vccd1
+ vccd1 net528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_1__f_wb_clk_i_X clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold61 team_10_WB.instance_to_wrap.gamelogic.red vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_10_WB.instance_to_wrap.host_row1\[46\] vssd1 vssd1 vccd1 vccd1 net550
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4118__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4268__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2253__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2690_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] _1336_ _1338_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4360_ clknet_leaf_11_wb_clk_i _0003_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3311_ net177 net552 vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_111_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4291_ clknet_leaf_16_wb_clk_i _0681_ _0280_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ net502 _1610_ net296 vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__a21oi_1
X_3173_ _0903_ _1298_ _1598_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_175_Right_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2124_ net211 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0927_ sky130_fd_sc_hd__mux2_1
XANTENNA__2428__B _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2055_ team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] net109 net135 team_10_WB.instance_to_wrap.dispFSM.guesses\[65\]
+ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_37_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2957_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] _0833_ net162 vssd1 vssd1 vccd1
+ vccd1 _1480_ sky130_fd_sc_hd__a41o_1
XFILLER_0_84_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1908_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1 vssd1 vccd1 vccd1
+ _0831_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2888_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] vssd1 vssd1 vccd1 vccd1
+ _1469_ sky130_fd_sc_hd__and3b_1
XANTENNA__2981__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4627_ net395 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
X_4494__305 vssd1 vssd1 vccd1 vccd1 _4494__305/HI net305 sky130_fd_sc_hd__conb_1
X_4558_ net369 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4489_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[46\]
+ _0472_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\]
+ sky130_fd_sc_hd__dfstp_1
X_3509_ net238 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__inv_2
X_4535__346 vssd1 vssd1 vccd1 vccd1 _4535__346/HI net346 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4410__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_0_170_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4090__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3860_ net273 vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2811_ _1413_ _1415_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__nor2_1
X_3791_ net279 vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2742_ team_10_WB.instance_to_wrap.clock_div.count\[15\] _1364_ _1366_ _1177_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[15\] sky130_fd_sc_hd__o211a_1
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2673_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ _1324_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__and3_1
X_4412_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[9\]
+ _0395_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_169_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4343_ clknet_leaf_22_wb_clk_i _0733_ _0332_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[66\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_185_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4274_ clknet_leaf_2_wb_clk_i _0664_ _0263_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3225_ net172 _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4433__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3156_ _1569_ _1574_ _1573_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__a21bo_1
X_3087_ _0790_ net206 vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__nor2_1
X_2107_ team_10_WB.instance_to_wrap.dispFSM.guesses\[13\] net144 net108 net530 vssd1
+ vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout267_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2038_ team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] net111 net137 team_10_WB.instance_to_wrap.dispFSM.msg\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[26\]
+ _0057_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout222_X net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3950__CLK clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1996__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3908__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4306__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3370__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4456__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3010_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\] net186 _1499_ net205
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[41\] sky130_fd_sc_hd__o211a_1
XFILLER_0_171_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3912_ net268 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1987__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3843_ net247 vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3774_ net293 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__inv_2
XANTENNA__3029__S net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2725_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ team_10_WB.instance_to_wrap.clock_div.count\[9\] _1351_ vssd1 vssd1 vccd1 vccd1
+ _1356_ sky130_fd_sc_hd__and4_2
XFILLER_0_124_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2656_ _1307_ _1316_ _1314_ _1228_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[1\]
+ sky130_fd_sc_hd__a211o_1
XANTENNA__2164__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2587_ net5 _0902_ _0904_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3361__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout115 net116 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_2
XFILLER_0_129_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4326_ clknet_leaf_17_wb_clk_i _0716_ _0315_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[49\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout126 _1191_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_4
Xfanout137 net142 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_2
Xfanout148 net150 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_4
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_4257_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[0\]
+ _0246_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3208_ net172 _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__nor2_1
X_4188_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[50\]
+ _0177_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[50\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2467__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3139_ _1286_ _1554_ _1565_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_107_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3973__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1978__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1978__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4329__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2927__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4479__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] vssd1 vssd1 vccd1 vccd1
+ net636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3352__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\] vssd1 vssd1 vccd1
+ vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2510_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net223 vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__and3_1
X_3490_ net248 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__inv_2
X_2441_ net504 net132 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\]
+ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__a22o_1
XANTENNA__3343__B1 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2372_ _1131_ _1135_ _1096_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__a21oi_1
X_4111_ clknet_leaf_9_wb_clk_i _0582_ _0110_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_4042_ clknet_leaf_14_wb_clk_i _0527_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3996__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3548__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout132_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3826_ net273 vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_15_wb_clk_i_X clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3757_ net278 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2708_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ net718 vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2385__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3688_ net236 vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2639_ _0946_ _1304_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[0\]
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4309_ clknet_leaf_14_wb_clk_i _0699_ _0298_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_58_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4151__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3325__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2256__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload8_A clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2990_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] net165 _1491_ net213
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[28\]
+ sky130_fd_sc_hd__o22a_1
X_1941_ net228 _0848_ _0851_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__o21ai_1
X_4660_ net428 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1872_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1 vccd1
+ _0797_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3611_ net260 vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4591_ net454 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2367__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3542_ net235 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__inv_2
X_3473_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] net169 _1844_ _1845_ vssd1 vssd1
+ vccd1 vccd1 _1846_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2424_ net197 _0942_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__nor2_4
X_2355_ _1128_ _1129_ _1126_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_4_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2286_ _0940_ _1064_ _1065_ _1063_ team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__a32o_1
X_4025_ clknet_leaf_33_wb_clk_i net558 _0072_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4174__CLK clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3809_ net284 vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4170__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4690__437 vssd1 vssd1 vccd1 vccd1 _4690__437/HI net437 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_189_Right_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3741__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2046__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3916__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4047__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3010__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4197__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2140_ _0822_ team_10_WB.instance_to_wrap.gamelogic.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0935_ sky130_fd_sc_hd__nand2_1
X_2071_ team_10_WB.instance_to_wrap.dispFSM.guesses\[41\] net110 net135 net696 vssd1
+ vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4255__Q team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2973_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] net126 _1486_ _1487_
+ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__nand4_4
X_1924_ net299 net3 vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__and2b_1
XFILLER_0_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4643_ net411 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4574_ net200 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3525_ net232 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_151_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3456_ team_10_WB.instance_to_wrap.host_row1\[46\] _1693_ net174 team_10_WB.instance_to_wrap.host_row2\[46\]
+ _1826_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3387_ team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] net167 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__a22o_1
X_2407_ _1168_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2338_ _0811_ _1093_ _1107_ _1108_ _1109_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_179_Left_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2269_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net212 vssd1 vssd1 vccd1
+ vccd1 _1051_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_162_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ clknet_leaf_21_wb_clk_i _0496_ net257 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_83_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_188_Left_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold40 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net496 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold51 team_10_WB.instance_to_wrap.host_row1\[64\] vssd1 vssd1 vccd1 vccd1 net507
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 net529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_10_WB.instance_to_wrap.host_row1\[57\] vssd1 vssd1 vccd1 vccd1 net518
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold95 team_10_WB.instance_to_wrap.host_row1\[66\] vssd1 vssd1 vccd1 vccd1 net551
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] vssd1 vssd1 vccd1
+ vccd1 net540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2518__C net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2990__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3310_ _1684_ _1689_ _1690_ net177 vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__or4b_1
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4290_ clknet_leaf_20_wb_clk_i net578 _0279_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_3241_ net468 _1642_ _1643_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__o21a_1
XFILLER_0_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3172_ _1290_ _1597_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] vssd1 vssd1 vccd1
+ vccd1 _1598_ sky130_fd_sc_hd__o21a_1
X_2123_ _0918_ _0925_ _0922_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_83_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2054_ team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] net111 net137 net653 vssd1
+ vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4641__409 vssd1 vssd1 vccd1 vccd1 _4641__409/HI net409 sky130_fd_sc_hd__conb_1
XANTENNA__4212__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3470__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2956_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\] net160 vssd1 vssd1 vccd1
+ vccd1 _1479_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1907_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] vssd1 vssd1 vccd1 vccd1
+ _0830_ sky130_fd_sc_hd__inv_2
X_2887_ _1222_ _1468_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[5\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_161_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4362__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout212_A team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4626_ net394 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_114_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4557_ net368 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3508_ net238 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__inv_2
X_4488_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[45\]
+ _0471_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_3439_ team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.dispFSM.guesses\[5\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2249__B1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3461__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput63 net200 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XANTENNA__2488__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4235__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3452__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2810_ _1415_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__inv_2
XANTENNA__4385__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3790_ net292 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2741_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2963__B2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3095__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4411_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[8\]
+ _0394_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_2672_ net528 _1324_ _1326_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4558__369 vssd1 vssd1 vccd1 vccd1 _4558__369/HI net369 sky130_fd_sc_hd__conb_1
X_4342_ clknet_leaf_18_wb_clk_i _0732_ _0331_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[65\]
+ sky130_fd_sc_hd__dfstp_1
X_4273_ clknet_leaf_0_wb_clk_i _0663_ _0262_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_185_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3224_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1632_ vssd1 vssd1 vccd1
+ vccd1 _1633_ sky130_fd_sc_hd__and2_1
.ends

