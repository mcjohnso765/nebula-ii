* NGSPICE file created from team_03.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

.subckt team_03 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XANTENNA__06990__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05903_ core.register_file.registers_state\[559\] core.register_file.registers_state\[527\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__mux2_1
XANTENNA__09523__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06883_ core.register_file.registers_state\[302\] core.register_file.registers_state\[270\]
+ core.register_file.registers_state\[430\] core.register_file.registers_state\[398\]
+ net847 net1076 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__mux4_1
X_09671_ _04845_ net286 net282 net1798 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__a22o_1
XANTENNA__08731__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ _04028_ _04064_ _04268_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__or4_1
X_05834_ core.register_file.registers_state\[784\] core.register_file.registers_state\[816\]
+ net697 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__mux2_1
XANTENNA__05832__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08553_ core.pc.current_pc\[30\] _04335_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nand2_1
XANTENNA__09287__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05765_ core.register_file.registers_state\[19\] core.register_file.registers_state\[51\]
+ net697 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07504_ _03582_ _03607_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__nand2_1
X_08484_ _04565_ _04566_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05696_ net950 net764 core.register_file.registers_state\[533\] vssd1 vssd1 vccd1
+ vccd1 _01801_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05848__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07435_ _03538_ _03539_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nand2_1
XANTENNA__05848__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1071_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07366_ net1094 core.register_file.registers_state\[730\] core.register_file.registers_state\[762\]
+ net836 net818 vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__o221a_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06317_ _01506_ _02421_ _02387_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_21_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09105_ net2493 net363 net352 _04861_ vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07297_ _03397_ _03401_ _03147_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06273__A1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09036_ net613 net216 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__and2_2
X_06248_ _02350_ _02352_ net646 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XANTENNA__11578__Q core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 core.CPU_DAT_I\[3\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10357__A0 _05109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06179_ net1044 core.register_file.registers_state\[102\] net750 _02283_ vssd1 vssd1
+ vccd1 vccd1 _02284_ sky130_fd_sc_hd__a31o_1
Xhold351 core.register_file.registers_state\[158\] vssd1 vssd1 vccd1 vccd1 net1670
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 core.register_file.registers_state\[286\] vssd1 vssd1 vccd1 vccd1 net1681
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _00004_ vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07222__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 core.register_file.registers_state\[401\] vssd1 vssd1 vccd1 vccd1 net1703
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09762__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 core.register_file.registers_state\[257\] vssd1 vssd1 vccd1 vccd1 net1714
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net823 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_2
Xfanout831 net834 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11812__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ core.decoder.inst\[27\] net2134 net894 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
Xfanout842 net846 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_2
XFILLER_0_99_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout853 net855 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_4
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_2
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09514__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 _01457_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_2
Xfanout897 _01398_ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ net558 _04945_ net456 net266 net2193 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__a32o_1
Xhold1040 core.register_file.registers_state\[211\] vssd1 vssd1 vccd1 vccd1 net2359
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 core.register_file.registers_state\[146\] vssd1 vssd1 vccd1 vccd1 net2370
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net1317 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
Xhold1062 core.register_file.registers_state\[472\] vssd1 vssd1 vccd1 vccd1 net2381
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06838__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1073 core.register_file.registers_state\[787\] vssd1 vssd1 vccd1 vccd1 net2392
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__A _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1084 core.register_file.registers_state\[83\] vssd1 vssd1 vccd1 vccd1 net2403
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06733__C1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 core.register_file.registers_state\[194\] vssd1 vssd1 vccd1 vccd1 net2414
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07523__A _01550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ clknet_leaf_24_clk net35 net1183 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09278__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ clknet_leaf_37_clk _01266_ net1222 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07810__X _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10713_ clknet_leaf_68_clk _00225_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[185\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ clknet_leaf_71_clk net1518 net1270 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10644_ clknet_leaf_53_clk _00156_ net1304 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08789__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10575_ clknet_leaf_83_clk _00087_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08253__A2 _04350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08073__B _03231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06264__A1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10348__A0 _05100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_19_clk_X clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08801__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11127_ clknet_leaf_22_clk _00639_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[599\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09505__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ clknet_leaf_67_clk _00570_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[530\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08713__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ net594 _02015_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06724__C1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07433__A _03536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09269__A1 _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05550_ net1026 _01648_ _01649_ _01654_ net932 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__o311a_1
XFILLER_0_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05481_ core.register_file.registers_state\[284\] core.register_file.registers_state\[316\]
+ core.register_file.registers_state\[412\] core.register_file.registers_state\[444\]
+ net699 net1019 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07220_ _03319_ _03323_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08264__A _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07151_ core.register_file.registers_state\[996\] core.register_file.registers_state\[964\]
+ net853 vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06102_ core.decoder.inst\[28\] net734 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07082_ _03181_ _03186_ _01462_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06033_ net1036 core.register_file.registers_state\[363\] net747 vssd1 vssd1 vccd1
+ vccd1 _02138_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11835__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10339__A0 _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06007__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07204__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__RESET_B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07984_ _03895_ _04088_ net492 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__mux2_1
XANTENNA__06963__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ _04918_ net286 net274 net1688 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__a22o_1
X_06935_ _03031_ _03034_ _03039_ net767 vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout377_A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ _04752_ net292 net284 net2124 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__a22o_1
X_06866_ core.register_file.registers_state\[814\] core.register_file.registers_state\[782\]
+ core.register_file.registers_state\[942\] core.register_file.registers_state\[910\]
+ net855 net1079 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ _04096_ _04679_ _04109_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11215__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05817_ _01920_ _01921_ net1031 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__o21ai_1
X_06797_ _02900_ _02901_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__nand2_1
X_09585_ _04935_ net402 net300 net2390 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1286_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ _04607_ _04613_ _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__nand3_1
X_05748_ _01849_ _01852_ net634 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08873__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ core.pc.current_pc\[22\] _02717_ net574 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05679_ net948 core.register_file.registers_state\[949\] net763 vssd1 vssd1 vccd1
+ vccd1 _01784_ sky130_fd_sc_hd__or3_1
XANTENNA__07140__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout809_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06494__A1 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06393__S net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07418_ _03517_ _03522_ net779 vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08398_ core.pc.current_pc\[15\] _04489_ net598 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__mux2_1
XANTENNA__08619__D_N _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_93_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ net1094 core.register_file.registers_state\[474\] core.register_file.registers_state\[506\]
+ net835 net1071 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__o221a_1
XANTENNA__08235__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10360_ _05112_ net1467 net235 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__mux2_1
XANTENNA__05310__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10042__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08902__A _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09019_ net742 net615 net206 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10291_ net14 net902 net796 net2282 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08621__B _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11481__SET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 _01224_ vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09735__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 _01229_ vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07746__A1 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 net164 vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__B1 _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05757__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_31_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 _01516_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_4
XANTENNA__09292__X _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout661 net663 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout672 net680 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_2
XFILLER_0_137_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08349__A _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08171__A1 _03890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11814_ clknet_leaf_72_clk _01315_ net1271 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09120__A0 _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11745_ clknet_leaf_35_clk _01257_ net1220 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11676_ clknet_leaf_35_clk _01188_ net1220 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10732__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11858__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10627_ clknet_leaf_73_clk _00139_ net1272 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_104_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06316__B _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06237__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10033__A2 _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10558_ clknet_leaf_96_clk _00070_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05996__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10489_ net1457 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09187__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10882__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09726__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05748__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07832__S1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06945__C1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06720_ net1108 core.register_file.registers_state\[338\] core.register_file.registers_state\[370\]
+ net858 net984 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06651_ core.register_file.registers_state\[532\] core.register_file.registers_state\[564\]
+ net889 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
X_05602_ net584 net593 _01665_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__or3_1
XANTENNA__11388__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06582_ _01866_ _02531_ net537 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__o21a_1
X_09370_ net2034 net330 net325 _04737_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05920__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09111__A0 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08321_ _04408_ _04412_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__nor2_1
X_05533_ net1035 core.register_file.registers_state\[218\] vssd1 vssd1 vccd1 vccd1
+ _01638_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07122__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ _04354_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__nor2_1
X_05464_ core.register_file.registers_state\[157\] net677 net641 _01568_ vssd1 vssd1
+ vccd1 vccd1 _01569_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07203_ core.register_file.registers_state\[2\] net884 net812 _03307_ vssd1 vssd1
+ vccd1 vccd1 _03308_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05411__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _02876_ _02902_ _03410_ _02875_ _02847_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__a311o_1
X_05395_ net1003 _01499_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__or2_2
XANTENNA__09414__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10029__A _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07134_ net994 core.register_file.registers_state\[68\] net884 core.register_file.registers_state\[100\]
+ net827 vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a221o_1
XANTENNA__10024__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06941__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11407__RESET_B net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ net992 core.register_file.registers_state\[583\] net879 core.register_file.registers_state\[615\]
+ net825 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09178__A0 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06016_ core.register_file.registers_state\[747\] core.register_file.registers_state\[715\]
+ net668 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XANTENNA__09717__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout494_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07625__X _03730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07967_ _03992_ _04025_ _04071_ _03688_ _04070_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout661_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout759_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _04893_ net2541 net278 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
X_06918_ net772 _03010_ _03021_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a22o_4
XFILLER_0_138_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06388__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ _03685_ _03994_ _04000_ _04001_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09350__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ net1001 _05011_ net460 net393 net2027 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__a32o_1
X_06849_ core.register_file.registers_state\[559\] core.register_file.registers_state\[527\]
+ net853 vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__mux2_1
XANTENNA__06164__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10211__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__S net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09568_ _04901_ net399 net301 net1991 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__a22o_1
XANTENNA__09102__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08519_ _04588_ _04599_ _04598_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10755__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07113__C1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ _04711_ net457 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06467__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07520__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ clknet_leaf_110_clk _01042_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1002\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_25_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06417__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05321__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11461_ clknet_leaf_101_clk _00973_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[933\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_34_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10412_ net1320 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_115_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11392_ clknet_leaf_57_clk _00904_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[864\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08632__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07967__B2 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07519__Y _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ _02343_ net1579 net233 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09169__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07248__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A gpio_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ net27 net904 net797 core.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11766__Q core.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07719__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06927__C1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07682__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__X _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_2
Xfanout491 _02487_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08144__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06155__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08807__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09402__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11728_ clknet_leaf_47_clk _01240_ net1291 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ clknet_leaf_47_clk _01171_ net1291 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05681__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold906 core.register_file.registers_state\[326\] vssd1 vssd1 vccd1 vccd1 net2225
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold917 core.register_file.registers_state\[642\] vssd1 vssd1 vccd1 vccd1 net2236
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 core.register_file.registers_state\[69\] vssd1 vssd1 vccd1 vccd1 net2247
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold939 core.register_file.registers_state\[628\] vssd1 vssd1 vccd1 vccd1 net2258
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07158__A _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_59_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11060__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08870_ _04891_ net2018 net373 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07821_ _03821_ _03925_ net481 vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09580__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07752_ _03717_ _03728_ net476 vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__mux2_1
XANTENNA__09332__A0 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05406__A core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06703_ net971 _02804_ _02807_ net776 vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a211o_1
X_07683_ _03781_ _03787_ net492 vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__mux2_1
XANTENNA__06146__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09883__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10031__B _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09422_ net2526 net205 net405 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
X_06634_ net826 _02735_ _02734_ net787 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__o211ai_1
XANTENNA__08717__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09353_ _05004_ net420 net414 net1742 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06565_ net1094 core.register_file.registers_state\[727\] core.register_file.registers_state\[759\]
+ net835 net818 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout242_A _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08304_ core.pc.current_pc\[6\] _04374_ core.pc.current_pc\[7\] vssd1 vssd1 vccd1
+ vccd1 _04404_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05516_ _01620_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06496_ _01632_ _01709_ _02600_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__o21ai_2
X_09284_ net2418 net212 net335 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05657__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08235_ _03319_ net577 _04337_ _02455_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05447_ net555 _01551_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1151_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1249_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08166_ _03685_ _04230_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__nand2_1
X_05378_ net971 _01481_ _01482_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07117_ net990 core.register_file.registers_state\[69\] net876 core.register_file.registers_state\[101\]
+ net824 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a221o_1
X_08097_ net513 _03872_ _04201_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload90 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_100_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07048_ net990 core.register_file.registers_state\[199\] net876 core.register_file.registers_state\[231\]
+ net809 vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a221o_1
XANTENNA__06621__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08602__D _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__Q core.IO_mod.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__C1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06385__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ net2298 net428 _04972_ net433 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09323__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05316__A core.decoder.inst\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10961_ clknet_leaf_74_clk _00473_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[433\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__A2 _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07334__C1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10892_ clknet_leaf_101_clk _00404_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[364\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06783__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05896__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05360__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10368__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05360__B2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06147__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05648__C1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11329__RESET_B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ clknet_leaf_60_clk _01025_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[985\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08633__Y _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11444_ clknet_leaf_56_clk _00956_ net1294 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[916\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08362__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11083__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11375_ clknet_leaf_79_clk _00887_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06612__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10326_ _05111_ net1598 net237 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05966__A3 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__Y _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10257_ net91 net914 vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__and2_1
XANTENNA__10964__RESET_B net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1220 net1224 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09562__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1231 net1232 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_4
X_10188_ net116 net918 net908 net1488 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a22o_1
Xfanout1242 net1250 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
Xfanout1253 net1278 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09624__C net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1264 net1268 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1275 net1276 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__clkbuf_4
Xfanout1286 net1313 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__buf_4
Xfanout1297 net1305 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_117_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09314__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08668__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09865__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05660__S net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05887__C1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08256__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06350_ net1122 _01409_ _01411_ net1015 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a22o_4
XANTENNA__06057__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05301_ core.decoder.inst\[30\] _01413_ _01414_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_44_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06281_ net1116 _01409_ _01411_ net1005 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a22o_4
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06300__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _02241_ _03139_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__nand2_1
XANTENNA__05654__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold703 core.register_file.registers_state\[357\] vssd1 vssd1 vccd1 vccd1 net2022
+ sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap411 _05057_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold714 core.register_file.registers_state\[248\] vssd1 vssd1 vccd1 vccd1 net2033
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09250__C1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold725 core.register_file.registers_state\[725\] vssd1 vssd1 vccd1 vccd1 net2044
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 core.ADR_I\[6\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06603__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold747 core.register_file.registers_state\[756\] vssd1 vssd1 vccd1 vccd1 net2066
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold758 core.register_file.registers_state\[677\] vssd1 vssd1 vccd1 vccd1 net2077
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09971_ net1471 core.CPU_DAT_O\[27\] net798 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__mux2_1
XANTENNA__07800__B1 _03902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold769 core.register_file.registers_state\[380\] vssd1 vssd1 vccd1 vccd1 net2088
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06603__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05811__C1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08922_ net2105 net367 _04921_ net431 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09553__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ _04887_ net2458 net372 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__mux2_1
XANTENNA__06367__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07804_ _03906_ _03907_ net494 vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__mux2_2
X_08784_ core.IO_mod.input_reg\[23\] net252 vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__nand2_1
XANTENNA__08108__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05996_ _02098_ _02100_ net622 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a21o_1
XANTENNA__09305__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ _03815_ _03816_ _03838_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout457_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ _03765_ _03770_ net494 vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_2
XFILLER_0_36_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09405_ net1900 _04885_ net405 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__mux2_1
X_06617_ net1105 core.register_file.registers_state\[725\] core.register_file.registers_state\[757\]
+ net851 net826 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__o221a_1
X_07597_ net500 _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout624_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05893__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ net1118 _04970_ net414 net1610 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06548_ net993 core.register_file.registers_state\[700\] net881 core.register_file.registers_state\[668\]
+ net825 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__o221a_1
XANTENNA__08734__X _04794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09084__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07095__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ net2195 _04886_ net337 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06479_ net1035 core.register_file.registers_state\[56\] net747 vssd1 vssd1 vccd1
+ vccd1 _02584_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _03840_ _03862_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06842__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09198_ _05001_ net360 net426 net1812 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout993_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ net265 _04251_ _04252_ _04253_ _04250_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__a311o_1
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06414__B net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09792__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11160_ clknet_leaf_5_clk _00672_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[632\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ _03917_ net588 vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nand2_1
XANTENNA__10943__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11091_ clknet_leaf_11_clk _00603_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[563\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10042_ net1481 net541 net520 _05121_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__a22o_1
XANTENNA__08898__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 core.register_file.registers_state\[953\] vssd1 vssd1 vccd1 vccd1 net1349
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold41 core.register_file.registers_state\[970\] vssd1 vssd1 vccd1 vccd1 net1360
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold52 core.register_file.registers_state\[1003\] vssd1 vssd1 vccd1 vccd1 net1371
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 core.register_file.registers_state\[993\] vssd1 vssd1 vccd1 vccd1 net1382
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 core.register_file.registers_state\[1000\] vssd1 vssd1 vccd1 vccd1 net1393
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 core.register_file.registers_state\[979\] vssd1 vssd1 vccd1 vccd1 net1404
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold96 core.register_file.registers_state\[1011\] vssd1 vssd1 vccd1 vccd1 net1415
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05581__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ clknet_leaf_55_clk _00456_ net1301 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[416\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08357__A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10875_ clknet_leaf_25_clk _00387_ net1191 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07086__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ clknet_leaf_66_clk _00939_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[899\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06046__C1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09783__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ clknet_leaf_93_clk _00870_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08820__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ net535 net1516 net236 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
X_11289_ clknet_leaf_55_clk _00801_ net1305 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[761\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09535__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05508__X _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09127__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08889__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 net1053 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1065 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__buf_2
Xfanout1072 core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
X_05850_ net631 _01951_ _01954_ net721 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a31o_1
Xfanout1083 net1090 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_33_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1094 net1096 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_2
X_05781_ net620 _01885_ _01884_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07520_ _03619_ net548 _03623_ _03616_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or4b_1
XFILLER_0_18_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07451_ core.register_file.registers_state\[607\] core.register_file.registers_state\[639\]
+ net700 vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06402_ _02503_ _02506_ net629 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__o21a_1
XANTENNA__10816__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07382_ core.register_file.registers_state\[25\] core.register_file.registers_state\[57\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__mux2_1
XANTENNA__09066__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09121_ _04889_ net2527 net347 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06333_ net955 core.register_file.registers_state\[32\] net765 vssd1 vssd1 vccd1
+ vccd1 _02438_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06264_ net953 core.register_file.registers_state\[68\] net710 core.register_file.registers_state\[100\]
+ net661 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a221o_1
XANTENNA__06824__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ net2372 net427 _05007_ net432 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08003_ _03658_ _03867_ _04104_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o211ai_4
X_06195_ net940 core.register_file.registers_state\[966\] vssd1 vssd1 vccd1 vccd1
+ _02300_ sky130_fd_sc_hd__and2_1
Xhold500 core.register_file.registers_state\[877\] vssd1 vssd1 vccd1 vccd1 net1819
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10037__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold511 core.register_file.registers_state\[526\] vssd1 vssd1 vccd1 vccd1 net1830
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 core.register_file.registers_state\[898\] vssd1 vssd1 vccd1 vccd1 net1841
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06037__C1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold533 core.register_file.registers_state\[910\] vssd1 vssd1 vccd1 vccd1 net1852
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09774__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 core.register_file.registers_state\[867\] vssd1 vssd1 vccd1 vccd1 net1863
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08730__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold555 core.register_file.registers_state\[557\] vssd1 vssd1 vccd1 vccd1 net1874
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 core.register_file.registers_state\[455\] vssd1 vssd1 vccd1 vccd1 net1885
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 core.register_file.registers_state\[852\] vssd1 vssd1 vccd1 vccd1 net1896
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 core.register_file.registers_state\[144\] vssd1 vssd1 vccd1 vccd1 net1907
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09954_ net1603 core.CPU_DAT_O\[10\] net801 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold599 core.register_file.registers_state\[872\] vssd1 vssd1 vccd1 vccd1 net1918
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09526__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08905_ _04746_ net736 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__and2_1
XANTENNA__10136__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ _04974_ net385 net378 net1748 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout574_A _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1200 core.register_file.registers_state\[643\] vssd1 vssd1 vccd1 vccd1 net2519
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 core.pc.current_pc\[1\] vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07001__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08836_ net731 _04878_ _04879_ net526 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__o211a_2
Xhold1222 core.register_file.registers_state\[730\] vssd1 vssd1 vccd1 vccd1 net2541
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06435__S0 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1233 core.register_file.registers_state\[731\] vssd1 vssd1 vccd1 vccd1 net2552
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ net571 net609 net214 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__and3_2
X_05979_ _02053_ _02083_ net585 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout839_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07718_ net476 _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08698_ _04670_ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__nor2_1
XANTENNA__11603__RESET_B net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07649_ net506 _03703_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06512__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05313__B _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10660_ clknet_leaf_77_clk _00172_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11741__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08905__A _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09319_ net558 _04945_ _05050_ net331 net2509 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ clknet_leaf_94_clk _00103_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06815__B2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout996_X net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06028__C1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11212_ clknet_leaf_103_clk _00724_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[684\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09765__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07240__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ clknet_leaf_65_clk _00655_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[615\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09780__A3 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__09517__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
X_11074_ clknet_leaf_78_clk _00586_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[546\]
+ sky130_fd_sc_hd__dfrtp_1
X_10025_ net594 _01745_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__nor2_4
XFILLER_0_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09296__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05504__A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10927_ clknet_leaf_83_clk _00439_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[399\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10858_ clknet_leaf_111_clk _00370_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[330\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09410__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07059__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_105_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10789_ clknet_leaf_87_clk _00301_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[261\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10063__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05609__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09756__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09220__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07231__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_4
XANTENNA__09508__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06070__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _03052_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__xor2_2
XANTENNA__05793__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05793__B2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05902_ core.register_file.registers_state\[815\] core.register_file.registers_state\[783\]
+ core.register_file.registers_state\[943\] core.register_file.registers_state\[911\]
+ net686 net1020 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09670_ _04839_ net287 net282 net2279 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__a22o_1
X_06882_ net794 _02985_ _02986_ _02984_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08731__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ _04074_ _04096_ _04679_ _04109_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__or4b_1
X_05833_ net1045 core.register_file.registers_state\[976\] core.register_file.registers_state\[1008\]
+ net673 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ _04626_ _04629_ core.pc.current_pc\[29\] net595 vssd1 vssd1 vccd1 vccd1 _00037_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06069__X _02174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05764_ net1047 core.register_file.registers_state\[179\] net674 core.register_file.registers_state\[147\]
+ net639 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a221o_1
XANTENNA__11764__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07105__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07503_ _03582_ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__or2_1
X_08483_ _01747_ _04552_ _04556_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05695_ net1055 core.register_file.registers_state\[565\] net756 vssd1 vssd1 vccd1
+ vccd1 _01800_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11014__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07434_ _03536_ _03537_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08725__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07365_ net803 _03468_ _03469_ net1082 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout322_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1064_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10054__B1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ net2285 net363 net352 _04856_ vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06316_ _02403_ _02420_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__nand2_4
XFILLER_0_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07296_ _03115_ _03143_ _03399_ _03087_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__and4b_1
XFILLER_0_115_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09035_ net2421 net429 _04996_ net1000 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06247_ net1059 core.register_file.registers_state\[612\] net754 _02351_ vssd1 vssd1
+ vccd1 vccd1 _02352_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1231_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07775__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07628__X _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09747__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold330 core.register_file.registers_state\[790\] vssd1 vssd1 vccd1 vccd1 net1649
+ sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ net940 core.register_file.registers_state\[70\] vssd1 vssd1 vccd1 vccd1 _02283_
+ sky130_fd_sc_hd__and2_1
Xhold341 _01204_ vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 core.register_file.registers_state\[550\] vssd1 vssd1 vccd1 vccd1 net1671
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 net157 vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold374 core.register_file.registers_state\[296\] vssd1 vssd1 vccd1 vccd1 net1693
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 core.register_file.registers_state\[822\] vssd1 vssd1 vccd1 vccd1 net1704
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 core.register_file.registers_state\[798\] vssd1 vssd1 vccd1 vccd1 net1715
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1117_X net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout810 net811 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout821 net823 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_4
X_09937_ core.decoder.inst\[26\] core.CPU_DAT_O\[26\] net893 vssd1 vssd1 vccd1 vccd1
+ _01090_ sky130_fd_sc_hd__mux2_1
XANTENNA__08970__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout832 net834 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_4
Xfanout843 net846 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout865 net874 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_4
Xfanout876 net882 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_4
X_09868_ _04943_ net388 net267 net1705 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__a22o_1
Xfanout887 net888 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__buf_4
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_4
Xhold1030 core.register_file.registers_state\[207\] vssd1 vssd1 vccd1 vccd1 net2349
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 core.register_file.registers_state\[149\] vssd1 vssd1 vccd1 vccd1 net2360
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1052 core.register_file.registers_state\[76\] vssd1 vssd1 vccd1 vccd1 net2371
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ net606 net210 vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__and2_1
XANTENNA__07081__S0 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1063 core.register_file.registers_state\[691\] vssd1 vssd1 vccd1 vccd1 net2382
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ net559 _04817_ net457 net270 net1646 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__a32o_1
Xhold1074 core.register_file.registers_state\[119\] vssd1 vssd1 vccd1 vccd1 net2393
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 core.register_file.registers_state\[461\] vssd1 vssd1 vccd1 vccd1 net2404
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ clknet_leaf_53_clk _01331_ net1300 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dfrtp_1
Xhold1096 core.register_file.registers_state\[907\] vssd1 vssd1 vccd1 vccd1 net2415
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07523__B _01709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ clknet_leaf_31_clk _00006_ net1201 vssd1 vssd1 vccd1 vccd1 core.ru.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08486__B1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10293__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10712_ clknet_leaf_3_clk _00224_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[184\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11692_ clknet_leaf_72_clk net1660 net1270 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08635__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10643_ clknet_leaf_12_clk _00155_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08789__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10574_ clknet_leaf_89_clk _00086_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07461__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05994__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09738__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09202__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10511__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08801__C net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11126_ clknet_leaf_61_clk _00638_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[598\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08961__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05775__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06972__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ clknet_leaf_74_clk _00569_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[529\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08713__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09405__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ net2495 net542 net521 _05104_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__a22o_1
XANTENNA__09910__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09632__C net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10140__A _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10284__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05480_ _01584_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06764__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05521__X _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11167__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09977__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07150_ core.register_file.registers_state\[868\] core.register_file.registers_state\[836\]
+ net854 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09441__A2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06101_ net582 _02204_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07081_ _03182_ _03183_ _03185_ _03184_ net805 net790 vssd1 vssd1 vccd1 vccd1 _03186_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09729__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06660__C1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06032_ core.register_file.registers_state\[299\] core.register_file.registers_state\[267\]
+ core.register_file.registers_state\[427\] core.register_file.registers_state\[395\]
+ net667 net1008 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06071__Y _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A3 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07755__A2 _03856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05409__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08952__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ _04085_ _04087_ net482 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__mux2_1
XANTENNA__05766__A1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06963__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09722_ _04916_ net290 net275 net2198 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__a22o_1
X_06934_ net970 _03035_ _03038_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a21o_1
XANTENNA__08704__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11266__RESET_B net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _04747_ net289 net283 net1994 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__a22o_1
X_06865_ net992 core.register_file.registers_state\[846\] net878 core.register_file.registers_state\[878\]
+ net1076 vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08604_ _04123_ _04677_ _04678_ _04172_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05816_ net1060 core.register_file.registers_state\[466\] core.register_file.registers_state\[498\]
+ net690 net1022 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__o221a_1
XANTENNA__10050__A _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ _04933_ net402 net300 net2064 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__a22o_1
X_06796_ _01957_ _02811_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06191__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07911__X _04016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ _04605_ _04608_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__nand2_1
X_05747_ net619 _01850_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout537_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__SET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08466_ core.pc.current_pc\[21\] _04551_ net596 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07140__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05678_ net950 core.register_file.registers_state\[661\] vssd1 vssd1 vccd1 vccd1
+ _01783_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07417_ _03518_ _03519_ _03521_ _03520_ net789 net816 vssd1 vssd1 vccd1 vccd1 _03522_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07691__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06494__A2 _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ _04488_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout704_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1067_X net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07348_ net1094 core.register_file.registers_state\[346\] core.register_file.registers_state\[378\]
+ net835 net978 vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09432__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10209__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07279_ _03352_ _03353_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08640__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08902__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09018_ net615 _04780_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10290_ net12 net904 net797 core.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 _01287_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__A1 _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 core.CPU_DAT_I\[5\] vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 core.register_file.registers_state\[4\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 core.register_file.registers_state\[987\] vssd1 vssd1 vccd1 vccd1 net1501
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10684__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 core.CPU_DAT_I\[1\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05319__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net642 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout673 net676 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout684 net685 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_2
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06706__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06182__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11813_ clknet_leaf_52_clk _01314_ net1303 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08636__Y _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05989__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11744_ clknet_leaf_35_clk _01256_ net1219 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05341__X _01449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09671__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11675_ clknet_leaf_35_clk _01187_ net1219 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ clknet_leaf_78_clk _00138_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10571__RESET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ clknet_leaf_17_clk _00069_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05445__A0 _01508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06172__X _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06613__A _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10488_ net1348 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10135__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07198__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08934__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06945__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ clknet_leaf_87_clk _00621_ net1229 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06759__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05663__S net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ _02753_ _02754_ net793 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07370__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07731__X _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05601_ net628 _01694_ _01705_ net717 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05381__C1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06581_ net771 _02674_ _02685_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a21oi_2
X_08320_ core.pc.current_pc\[9\] _04413_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05532_ net938 core.register_file.registers_state\[250\] net757 vssd1 vssd1 vccd1
+ vccd1 _01637_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07122__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10557__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08251_ _02386_ _04353_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__nor2_1
XANTENNA__07610__C net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05463_ net1051 core.register_file.registers_state\[189\] vssd1 vssd1 vccd1 vccd1
+ _01568_ sky130_fd_sc_hd__and2_1
XANTENNA__08870__A0 _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11802__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07202_ core.register_file.registers_state\[34\] net856 vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05411__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ net527 _03986_ _04279_ _04285_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06881__C1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05394_ _01407_ _01417_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__or2_2
XANTENNA__10029__B _02560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload57_A clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07133_ core.register_file.registers_state\[36\] core.register_file.registers_state\[4\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__mux2_1
XANTENNA__06228__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_65_clk_X clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07064_ net992 core.register_file.registers_state\[711\] net878 core.register_file.registers_state\[743\]
+ net809 vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05987__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05987__B2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06015_ core.register_file.registers_state\[683\] core.register_file.registers_state\[651\]
+ net668 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1027_A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08925__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05739__B2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _04009_ _04013_ _04058_ _04011_ _02487_ net480 vssd1 vssd1 vccd1 vccd1 _04071_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_96_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ net211 net1961 net281 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
X_06917_ _01462_ _03015_ _03016_ net768 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ net507 _03640_ _03651_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout654_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09350__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09636_ net2056 net391 _05078_ net998 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__a22o_1
X_06848_ core.register_file.registers_state\[623\] core.register_file.registers_state\[591\]
+ net853 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06164__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ _04899_ net401 net300 net2024 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05911__A1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06779_ net1097 core.register_file.registers_state\[464\] core.register_file.registers_state\[496\]
+ net839 net1073 vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout919_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08518_ _04573_ _04578_ _04587_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__or3_1
XANTENNA__07113__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _04711_ net456 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__and2_1
XANTENNA__09653__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05602__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08449_ _04532_ _04534_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06417__B _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05675__B1 _01779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05321__B core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ clknet_leaf_81_clk _00972_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[932\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ net1344 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_115_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05690__A3 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ clknet_leaf_41_clk _00903_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08632__B net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ net535 net1531 net232 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05978__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10273_ net24 net904 net797 core.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08916__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A gpio_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout470 _05127_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout481 _02517_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 _02486_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08144__A2 _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06155__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07551__X _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08807__B _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10752__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06167__X _02272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05512__A _01395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11727_ clknet_leaf_47_clk _01239_ net1306 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10254__A3 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ clknet_leaf_46_clk _01170_ net1291 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10609_ clknet_leaf_72_clk _00121_ net1269 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11589_ clknet_leaf_28_clk _01101_ net1197 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold907 core.register_file.registers_state\[228\] vssd1 vssd1 vccd1 vccd1 net2226
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold918 core.register_file.registers_state\[184\] vssd1 vssd1 vccd1 vccd1 net2237
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 core.register_file.registers_state\[590\] vssd1 vssd1 vccd1 vccd1 net2248
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05969__B2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08907__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ net505 _03674_ _03672_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07186__A3 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10190__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _03700_ _03711_ _03724_ _03704_ net479 net491 vssd1 vssd1 vccd1 vccd1 _03856_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_100_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_92_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
X_06702_ _02805_ _02806_ net1085 vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__o21a_1
XANTENNA__05406__B net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ _03784_ _03786_ net482 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__mux2_1
XANTENNA__10031__C _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ net1921 net213 net407 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06633_ _02736_ _02737_ net794 vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_138_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05354__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09352_ net1120 _05002_ net415 net1764 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09096__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06564_ net804 _02667_ _02668_ net1090 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08303_ core.pc.current_pc\[6\] core.pc.current_pc\[7\] _04374_ vssd1 vssd1 vccd1
+ vccd1 _04403_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05515_ _01496_ _01618_ _01366_ _01418_ _01489_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__o2111a_2
XANTENNA__08843__A0 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ net2536 net205 net335 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__mux2_1
X_06495_ _02534_ _02599_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout235_A _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ _03319_ _04335_ _04338_ _02455_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05446_ core.decoder.inst\[29\] net898 net593 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__a21o_1
XANTENNA__06952__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08733__A core.IO_mod.input_reg\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05752__S0 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09399__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08165_ net528 _04269_ _03410_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__or3b_1
X_05377_ net1099 core.register_file.registers_state\[606\] core.register_file.registers_state\[638\]
+ net843 net805 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout402_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07116_ _03218_ _03220_ net785 vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08096_ net513 _04106_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_110_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload80 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__inv_8
XANTENNA_clkbuf_leaf_45_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload91 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__inv_12
X_07047_ net992 core.register_file.registers_state\[71\] net879 core.register_file.registers_state\[103\]
+ net825 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1311_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A1 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11210__RESET_B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__C1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06385__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net568 _04971_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__and2_1
XANTENNA__10181__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ net490 _04012_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nand2_1
XANTENNA__05593__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_108_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_103_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05316__B core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ clknet_leaf_108_clk _00472_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[432\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08908__A _04751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09874__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09619_ net2473 net394 _05071_ net1000 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__a22o_1
X_10891_ clknet_leaf_110_clk _00403_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[363\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05896__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09087__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10236__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ clknet_leaf_4_clk _01024_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[984\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08643__A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11443_ clknet_leaf_11_clk _00955_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[915\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11369__RESET_B net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11374_ clknet_leaf_90_clk _00886_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[846\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11777__Q core.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ _05110_ net183 net239 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
X_10256_ net1125 net1977 net910 _05236_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__a31o_1
Xfanout1210 net1213 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_4
Xfanout1221 net1223 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1232 net1236 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_2
X_10187_ net115 net918 net908 net1525 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a22o_1
Xfanout1243 net1246 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10172__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1254 net1257 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1265 net1267 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1276 net1277 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__clkbuf_2
Xfanout1287 net1313 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_58_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09314__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1298 net1301 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09413__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09640__C net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05887__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09078__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06338__A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05300_ _01413_ _01414_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__or2_1
XANTENNA__05639__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06280_ net586 net535 _02382_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_44_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold704 core.register_file.registers_state\[638\] vssd1 vssd1 vccd1 vccd1 net2023
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06073__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold715 core.register_file.registers_state\[420\] vssd1 vssd1 vccd1 vccd1 net2034
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08840__X _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold726 core.register_file.registers_state\[573\] vssd1 vssd1 vccd1 vccd1 net2045
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 core.register_file.registers_state\[664\] vssd1 vssd1 vccd1 vccd1 net2056
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09970_ net1553 core.CPU_DAT_O\[26\] net800 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__mux2_1
XANTENNA__07800__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07261__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold748 core.register_file.registers_state\[645\] vssd1 vssd1 vccd1 vccd1 net2067
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11039__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold759 core.register_file.registers_state\[809\] vssd1 vssd1 vccd1 vccd1 net2078
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08921_ net563 net222 net735 vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07013__C1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__D1 _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ net741 _04758_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06367__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__inv_2
XANTENNA__05417__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08783_ net732 _03985_ net526 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05575__C1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05995_ core.register_file.registers_state\[12\] net675 net655 _02099_ vssd1 vssd1
+ vccd1 vccd1 _02100_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_49_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
X_07734_ _03815_ _03816_ _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__o21a_2
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06119__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06119__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09856__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ net484 _03767_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__RESET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09404_ net2117 _04884_ net407 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1094_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06616_ net1105 core.register_file.registers_state\[597\] core.register_file.registers_state\[629\]
+ net851 net811 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__o221a_1
X_07596_ _02530_ _03140_ _03630_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__or3_4
XFILLER_0_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09608__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ net1118 _04968_ net414 net1985 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__a22o_1
XANTENNA__10218__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06547_ core.register_file.registers_state\[540\] core.register_file.registers_state\[572\]
+ net881 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout617_A _01524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1261_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ net2225 _04885_ net335 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06478_ net1035 core.register_file.registers_state\[184\] net666 core.register_file.registers_state\[152\]
+ net637 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08217_ _03946_ _04318_ _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05429_ _01530_ _01533_ _01522_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a21oi_1
X_09197_ _04999_ net354 net423 net2118 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08148_ _04084_ _04025_ _03950_ _03797_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07478__S0 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10217__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06055__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08079_ net495 _04183_ _04181_ _03688_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1314_X net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10110_ net1124 net556 vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11090_ clknet_leaf_67_clk _00602_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[562\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11670__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _03566_ _03580_ net594 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_41_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold20 core.register_file.registers_state\[947\] vssd1 vssd1 vccd1 vccd1 net1339
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 core.register_file.registers_state\[935\] vssd1 vssd1 vccd1 vccd1 net1350
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold42 core.register_file.registers_state\[941\] vssd1 vssd1 vccd1 vccd1 net1361
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold53 core.register_file.registers_state\[22\] vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 core.register_file.registers_state\[1010\] vssd1 vssd1 vccd1 vccd1 net1383
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05566__C1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold75 core.register_file.registers_state\[960\] vssd1 vssd1 vccd1 vccd1 net1394
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 core.register_file.registers_state\[21\] vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 core.register_file.registers_state\[972\] vssd1 vssd1 vccd1 vccd1 net1416
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09847__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943_ clknet_leaf_14_clk _00455_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[415\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06429__Y _02534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05869__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_10874_ clknet_leaf_5_clk _00386_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[346\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09480__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07491__C1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11426_ clknet_leaf_79_clk _00938_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[898\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09232__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ clknet_leaf_20_clk _00869_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[829\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08820__B net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09408__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ _02421_ net1543 net236 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11288_ clknet_leaf_5_clk _00800_ net1146 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[760\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09635__C net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10239_ net81 net921 vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__and2_1
XANTENNA__06349__A1 _01506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1051 net1052 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
Xfanout1062 net1065 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05557__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_4
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_8
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09299__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__S net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05780_ core.register_file.registers_state\[531\] core.register_file.registers_state\[563\]
+ core.register_file.registers_state\[659\] core.register_file.registers_state\[691\]
+ net697 net654 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux4_1
XANTENNA__08548__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07450_ core.register_file.registers_state\[543\] core.register_file.registers_state\[575\]
+ net700 vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06521__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06521__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06401_ net625 _02504_ _02505_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07381_ net1089 _03482_ _03485_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__o21ai_1
X_09120_ _04888_ net2267 net347 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06332_ net1063 core.register_file.registers_state\[128\] net691 core.register_file.registers_state\[160\]
+ net663 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09471__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09051_ net565 net603 net205 vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__and3_1
X_06263_ _02365_ _02367_ net619 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08002_ _03872_ _04018_ _04025_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_5_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06194_ net1045 core.register_file.registers_state\[870\] net750 _02298_ vssd1 vssd1
+ vccd1 vccd1 _02299_ sky130_fd_sc_hd__a31o_1
XANTENNA__09223__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold501 core.register_file.registers_state\[760\] vssd1 vssd1 vccd1 vccd1 net1820
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10037__B _01582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold512 core.register_file.registers_state\[683\] vssd1 vssd1 vccd1 vccd1 net1831
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold523 core.register_file.registers_state\[446\] vssd1 vssd1 vccd1 vccd1 net1842
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11693__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold534 core.register_file.registers_state\[441\] vssd1 vssd1 vccd1 vccd1 net1853
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 core.register_file.registers_state\[736\] vssd1 vssd1 vccd1 vccd1 net1864
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 core.IO_mod.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06588__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06588__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08730__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 core.register_file.registers_state\[829\] vssd1 vssd1 vccd1 vccd1 net1886
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07627__A _03697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold578 core.register_file.registers_state\[435\] vssd1 vssd1 vccd1 vccd1 net1897
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net2090 net2068 net798 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
Xhold589 core.register_file.registers_state\[535\] vssd1 vssd1 vccd1 vccd1 net1908
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09526__A1 _04851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ net2451 net369 _04909_ net436 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__a22o_1
XANTENNA__10053__A _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09884_ _04972_ net390 net377 net1899 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1107_A core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 core.register_file.registers_state\[311\] vssd1 vssd1 vccd1 vccd1 net2520
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 core.register_file.registers_state\[59\] vssd1 vssd1 vccd1 vccd1 net2531
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ net731 net255 vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05548__C1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06435__S1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1223 core.register_file.registers_state\[827\] vssd1 vssd1 vccd1 vccd1 net2542
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 core.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08729__Y _04790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ net609 net214 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05978_ net721 _02066_ _02075_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__o22a_4
XFILLER_0_135_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07717_ _03661_ _03662_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_101_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ net728 _04123_ net525 _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout734_A _01412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1097_X net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ net452 _03080_ net444 net501 vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ _02346_ _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__nand2_2
XANTENNA__08905__B net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09318_ core.register_file.registers_state\[375\] net474 net544 vssd1 vssd1 vccd1
+ vccd1 _05050_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10590_ clknet_leaf_92_clk _00102_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09462__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05610__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09249_ net558 _04862_ _05040_ net339 net2467 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08017__A1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09214__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ clknet_leaf_107_clk _00723_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[683\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07225__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06123__S0 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06579__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11142_ clknet_leaf_99_clk _00654_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[614\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__clkbuf_4
X_11073_ clknet_leaf_85_clk _00585_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[545\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
X_10024_ net1525 net542 net521 _05112_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__a22o_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05539__C1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06200__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ clknet_leaf_88_clk _00438_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[398\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06503__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06503__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10857_ clknet_leaf_38_clk _00369_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[329\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10788_ clknet_leaf_80_clk _00300_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[260\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09453__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10063__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06267__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09205__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08831__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07216__C1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11409_ clknet_leaf_66_clk _00921_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[881\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09138__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06351__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05778__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06950_ _02146_ _03054_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06990__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07734__X _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05901_ _02004_ _02005_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__and2_1
XANTENNA__11096__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06881_ net991 core.register_file.registers_state\[206\] net877 core.register_file.registers_state\[238\]
+ net808 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08620_ _03734_ _04694_ _03811_ _04692_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__or4b_1
X_05832_ core.register_file.registers_state\[912\] core.register_file.registers_state\[944\]
+ net697 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
XANTENNA__08731__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ net208 _04627_ _04628_ net595 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__o31a_1
X_05763_ core.decoder.inst\[19\] net896 _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_72_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07502_ net549 vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08482_ _01710_ _04564_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__or2_1
XANTENNA__09692__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05694_ net1055 core.register_file.registers_state\[693\] net764 _01783_ net928 vssd1
+ vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07433_ _03536_ _03537_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__nand2_1
XANTENNA__10933__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07364_ net987 core.register_file.registers_state\[698\] net868 core.register_file.registers_state\[666\]
+ net818 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__o221a_1
XANTENNA__09444__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09103_ net2378 net365 net360 _04850_ vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__a22o_1
X_06315_ _02419_ net718 _02412_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__or3b_4
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08798__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07295_ _03115_ _03143_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout315_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09034_ net743 net465 _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__and3_1
X_06246_ net951 core.register_file.registers_state\[580\] vssd1 vssd1 vccd1 vccd1
+ _02351_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06960__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold320 core.register_file.registers_state\[363\] vssd1 vssd1 vccd1 vccd1 net1639
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06177_ _02279_ _02281_ net617 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__o21ai_1
Xhold331 core.register_file.registers_state\[775\] vssd1 vssd1 vccd1 vccd1 net1650
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 core.register_file.registers_state\[925\] vssd1 vssd1 vccd1 vccd1 net1661
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1224_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 core.register_file.registers_state\[415\] vssd1 vssd1 vccd1 vccd1 net1672
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 core.register_file.registers_state\[908\] vssd1 vssd1 vccd1 vccd1 net1683
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06261__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold375 core.register_file.registers_state\[803\] vssd1 vssd1 vccd1 vccd1 net1694
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_4
Xhold386 core.register_file.registers_state\[886\] vssd1 vssd1 vccd1 vccd1 net1705
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold397 net181 vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _01460_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06430__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08970__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ core.decoder.inst\[25\] net1678 net891 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10109__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1012_X net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_4
Xfanout844 net846 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_2
Xfanout855 net861 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_4
Xfanout866 net868 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_4
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 net882 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
X_09867_ _04941_ net388 net267 net1972 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__a22o_1
Xhold1020 core.register_file.registers_state\[92\] vssd1 vssd1 vccd1 vccd1 net2339
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net890 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_4
Xfanout899 net901 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
Xhold1031 core.register_file.registers_state\[465\] vssd1 vssd1 vccd1 vccd1 net2350
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 core.register_file.registers_state\[244\] vssd1 vssd1 vccd1 vccd1 net2361
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ net732 _03964_ net526 _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__o211a_2
Xhold1053 core.register_file.registers_state\[151\] vssd1 vssd1 vccd1 vccd1 net2372
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07081__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1064 core.register_file.registers_state\[113\] vssd1 vssd1 vccd1 vccd1 net2383
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ _04812_ net388 net271 net2012 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__a22o_1
XANTENNA__06733__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1075 core.register_file.registers_state\[94\] vssd1 vssd1 vccd1 vccd1 net2394
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 core.register_file.registers_state\[345\] vssd1 vssd1 vccd1 vccd1 net2405
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 core.register_file.registers_state\[833\] vssd1 vssd1 vccd1 vccd1 net2416
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__C _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ net572 net608 net217 vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11760_ clknet_leaf_31_clk _00005_ net1201 vssd1 vssd1 vccd1 vccd1 core.ru.state\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09683__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10293__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ clknet_leaf_20_clk _00223_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11691_ clknet_leaf_71_clk net1541 net1270 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08635__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10642_ clknet_leaf_69_clk _00154_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09435__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08789__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10573_ clknet_leaf_106_clk _00085_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05486__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07267__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__B2 _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__Q core.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11125_ clknet_leaf_64_clk _00637_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[597\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08961__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07554__X _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_X net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ clknet_leaf_104_clk _00568_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[528\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _01502_ _02051_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__nor2_2
XANTENNA__08713__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__A _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06724__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06724__B2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05932__C1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09674__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09421__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10284__B2 core.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ clknet_leaf_18_clk _00421_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11889_ clknet_leaf_70_clk _01358_ net1276 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05250__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__B2 _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06100_ core.decoder.inst\[29\] net734 net582 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07080_ core.register_file.registers_state\[998\] core.register_file.registers_state\[966\]
+ net839 vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06031_ _02132_ _02135_ net628 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08952__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07982_ net504 _03645_ _03783_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__o21ai_1
XANTENNA__05409__B net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06963__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06933_ net1083 _03036_ _03037_ net775 vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__a31o_1
X_09721_ _04914_ net290 net274 net2063 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09901__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _04742_ net289 net283 net2077 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__a22o_1
X_06864_ net992 core.register_file.registers_state\[974\] net878 core.register_file.registers_state\[1006\]
+ net983 vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__a221o_1
X_08603_ _04139_ _04155_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05815_ net1061 core.register_file.registers_state\[338\] core.register_file.registers_state\[370\]
+ net691 net930 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__o221a_1
X_09583_ _04931_ net397 net299 net2069 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__a22o_1
XANTENNA__06020__S net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10050__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06795_ net768 _02899_ _02887_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__o21a_4
XANTENNA__05923__C1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08534_ _01584_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__xnor2_1
X_05746_ net1063 core.register_file.registers_state\[212\] core.register_file.registers_state\[244\]
+ net691 net662 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06955__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09665__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08736__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08465_ _04550_ _04542_ net231 vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__mux2_1
XANTENNA__10275__B2 core.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05677_ net1028 net899 net593 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout432_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07140__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07416_ core.register_file.registers_state\[920\] core.register_file.registers_state\[952\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11111__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ _04487_ _04480_ net230 vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__mux2_1
XANTENNA__07691__A2 _03791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__C _03412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ core.register_file.registers_state\[282\] core.register_file.registers_state\[314\]
+ core.register_file.registers_state\[410\] core.register_file.registers_state\[442\]
+ net868 net1069 vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06326__S0 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09432__A3 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07278_ net497 _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08640__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout899_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11261__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ core.register_file.registers_state\[139\] net427 _04984_ net998 vssd1 vssd1
+ vccd1 vccd1 _00179_ sky130_fd_sc_hd__a22o_1
X_06229_ net941 core.register_file.registers_state\[677\] core.register_file.registers_state\[645\]
+ net698 net655 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10870__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold150 net199 vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 _01206_ vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold172 net139 vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 net150 vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 _01202_ vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05319__B net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _01522_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout641 net642 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_4
X_09919_ core.decoder.inst\[8\] core.CPU_DAT_O\[8\] net892 vssd1 vssd1 vccd1 vccd1
+ _01072_ sky130_fd_sc_hd__mux2_1
Xfanout652 net653 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 net664 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_4
XANTENNA__08156__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 net675 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10979__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout685 _01514_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout696 net716 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11812_ clknet_leaf_71_clk _01313_ net1274 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08646__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09656__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11743_ clknet_leaf_35_clk _01255_ net1219 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11674_ clknet_leaf_35_clk _01186_ net1219 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10018__B2 _05109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07419__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10625_ clknet_leaf_86_clk _00137_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07696__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08092__C1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10556_ clknet_leaf_40_clk _00068_ net1218 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05445__A1 _01549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ net1379 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09187__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07198__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06945__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ clknet_leaf_74_clk _00620_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[580\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09416__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11520__SET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11039_ clknet_leaf_14_clk _00551_ net1177 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[511\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09895__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05600_ _01696_ _01699_ _01704_ net621 net631 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06580_ net779 _02679_ _02684_ net767 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__o211a_1
XANTENNA__09647__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05531_ net1034 core.register_file.registers_state\[90\] core.register_file.registers_state\[122\]
+ net670 net638 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07122__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08250_ _02386_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05462_ net1026 _01566_ net721 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07673__A2 _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06076__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07201_ net1111 core.register_file.registers_state\[130\] net856 core.register_file.registers_state\[162\]
+ net827 vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08181_ net527 _03986_ _04279_ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06881__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05393_ _01417_ _01425_ _01491_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__or3_4
XANTENNA__06308__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07132_ net1111 core.register_file.registers_state\[132\] net856 core.register_file.registers_state\[164\]
+ net827 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07063_ net824 _03166_ _03167_ net975 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__o211a_1
XANTENNA__06633__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput200 net200 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_101_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06014_ core.register_file.registers_state\[619\] core.register_file.registers_state\[587\]
+ net668 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
XANTENNA__06015__S net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08925__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10193__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _03854_ _04018_ _04067_ _04069_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_96_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ net212 net2543 net278 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
X_06916_ net974 _03017_ _03020_ net776 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a211o_1
X_07896_ _03798_ _03843_ _03858_ _03980_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09886__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ net742 _05008_ net456 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__and3_1
X_06847_ core.register_file.registers_state\[751\] core.register_file.registers_state\[719\]
+ net853 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1291_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06778_ net1097 core.register_file.registers_state\[336\] core.register_file.registers_state\[368\]
+ net833 net980 vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__o221a_1
XANTENNA__09638__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ net1121 net601 _05062_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05911__A2 _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ _04596_ _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05729_ net955 core.register_file.registers_state\[564\] net765 vssd1 vssd1 vccd1
+ vccd1 _01834_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07113__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ net544 net474 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__and2b_4
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_X net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05602__B net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ _04515_ _04533_ _04532_ _04524_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06467__A3 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__X _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06321__C1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06872__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08379_ _04470_ _04471_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05321__C core.decoder.inst\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10410_ net1337 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10651__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11777__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ clknet_leaf_95_clk _00902_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[862\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09810__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10341_ _02421_ net1511 net234 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09169__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10272_ net13 net905 net797 core.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11007__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08916__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10184__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 _05060_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_2
Xfanout471 _05127_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_2
Xfanout482 _02516_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout493 _02486_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09877__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__X _03937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08144__A3 _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06595__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05352__X _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09644__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ clknet_leaf_48_clk _01238_ net1306 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ clknet_leaf_47_clk _01169_ net1306 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ clknet_leaf_107_clk _00120_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11588_ clknet_leaf_26_clk _01100_ net1193 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09801__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09000__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold908 core.register_file.registers_state\[197\] vssd1 vssd1 vccd1 vccd1 net2227
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__A2 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10539_ clknet_leaf_109_clk _00051_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold919 core.register_file.registers_state\[178\] vssd1 vssd1 vccd1 vccd1 net2238
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08907__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06918__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10175__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05527__X _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09580__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07750_ _03687_ _03854_ _03852_ _03847_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a211o_1
XANTENNA__09868__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06701_ net1097 core.register_file.registers_state\[467\] core.register_file.registers_state\[499\]
+ net840 net1074 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__o221a_1
X_07681_ net507 _03641_ _03785_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06777__S0 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06632_ net1105 core.register_file.registers_state\[213\] core.register_file.registers_state\[245\]
+ net851 net826 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__o221a_1
X_09420_ net2201 _04891_ net407 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05354__B1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08286__A _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06551__C1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09351_ net1115 net463 _05000_ net413 net1537 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__a32o_1
X_06563_ net987 core.register_file.registers_state\[695\] net874 core.register_file.registers_state\[663\]
+ net818 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08302_ _04400_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__and2_1
X_05514_ _01496_ _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09282_ net2168 net213 net337 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
XANTENNA__10674__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06494_ _02561_ _02598_ net537 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08233_ _01380_ _04335_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05445_ _01508_ _01549_ net584 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout228_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05752__S1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _03403_ _03407_ _03409_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05376_ net1099 core.register_file.registers_state\[734\] core.register_file.registers_state\[766\]
+ net841 net819 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__o221a_1
XANTENNA__06534__A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07115_ core.register_file.registers_state\[5\] net870 net809 _03219_ vssd1 vssd1
+ vccd1 vccd1 _03220_ sky130_fd_sc_hd__o211a_1
X_08095_ _04017_ _04199_ _04198_ _04194_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__o211a_4
XANTENNA__10056__A _04215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1137_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload70 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_110_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ _03148_ _03150_ net786 vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload81 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload92 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_fanout597_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09020__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10166__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1304_A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__B2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout764_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ net611 _04741_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07948_ _04024_ _04049_ _04050_ _03621_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09323__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__RESET_B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05316__C core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _03686_ _03974_ _03982_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07334__A1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07371__Y _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08908__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ net743 _04989_ net459 vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10890_ clknet_leaf_111_clk _00402_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[362\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06709__A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05896__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09549_ net219 net2277 net304 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08924__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06147__C net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05648__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11511_ clknet_leaf_6_clk _01023_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[983\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05648__B2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08643__B _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11442_ clknet_leaf_64_clk _00954_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[914\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11373_ clknet_leaf_0_clk _00885_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[845\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08062__A2 _03201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input60_A gpio_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ _05109_ net1716 net238 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10255_ net89 net914 vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09011__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_4
Xfanout1211 net1213 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_2
Xfanout1222 net1223 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_4
X_10186_ net114 net918 net908 net1495 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a22o_1
Xfanout1233 net1235 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_4
Xfanout1244 net1246 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08770__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1255 net1257 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1266 net1267 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08658__X _04730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1277 net1278 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1288 net1292 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06781__C1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_4
Xfanout1299 net1301 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09865__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload6_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10697__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06533__C1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05887__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09078__B2 _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10902__RESET_B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05639__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ clknet_leaf_54_clk net1573 net1299 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06300__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08553__B _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08589__B1 _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold705 core.register_file.registers_state\[608\] vssd1 vssd1 vccd1 vccd1 net2024
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold716 core.register_file.registers_state\[303\] vssd1 vssd1 vccd1 vccd1 net2035
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold727 core.register_file.registers_state\[352\] vssd1 vssd1 vccd1 vccd1 net2046
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold738 core.register_file.registers_state\[366\] vssd1 vssd1 vccd1 vccd1 net2057
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold749 core.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__A2 _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05811__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ net222 net735 vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09002__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_X clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07185__A _03289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08210__C1 _04312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _04886_ net2259 net373 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__mux2_1
XANTENNA__07564__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11472__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07802_ _03746_ _03779_ net478 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
XANTENNA__11008__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05417__B net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05994_ net1049 core.register_file.registers_state\[44\] net750 vssd1 vssd1 vccd1
+ vccd1 _02099_ sky130_fd_sc_hd__and3_1
X_08782_ net2329 net468 net437 _04834_ vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09305__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ _03697_ _03820_ _03837_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_75_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10320__A0 _05105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ net478 _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__or2_1
XANTENNA__06529__A _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09403_ net2095 net223 net408 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06615_ _02717_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__nor2_1
X_07595_ _03698_ _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout345_A _05027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06546_ net1087 _02647_ _02650_ net1067 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__o211a_1
X_09334_ net1118 _04966_ net414 net1687 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10643__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09265_ net1990 _04884_ net337 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__mux2_1
X_06477_ net1025 _02574_ net721 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout512_A _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1254_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08216_ _03985_ _04317_ _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__nor3_1
X_05428_ net962 _01532_ _01531_ net927 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a211o_1
X_09196_ _04997_ net360 net426 net1662 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ net494 _04236_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05359_ net1098 core.register_file.registers_state\[94\] core.register_file.registers_state\[126\]
+ net842 net806 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__o221a_1
XANTENNA__08044__A2 _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_X net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07478__S1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ _04145_ _04182_ net479 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09792__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07029_ net1083 _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_8_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10040_ net1567 net542 net521 _05120_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11431__RESET_B net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10233__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 core.register_file.registers_state\[934\] vssd1 vssd1 vccd1 vccd1 net1329
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 core.register_file.registers_state\[977\] vssd1 vssd1 vccd1 vccd1 net1340
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 core.register_file.registers_state\[982\] vssd1 vssd1 vccd1 vccd1 net1351
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold43 core.register_file.registers_state\[1023\] vssd1 vssd1 vccd1 vccd1 net1362
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05566__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold54 core.register_file.registers_state\[1017\] vssd1 vssd1 vccd1 vccd1 net1373
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 core.register_file.registers_state\[940\] vssd1 vssd1 vccd1 vccd1 net1384
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold76 core.ADR_I\[8\] vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__A _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 core.register_file.registers_state\[13\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 core.register_file.registers_state\[983\] vssd1 vssd1 vccd1 vccd1 net1417
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08638__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10311__A0 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10942_ clknet_leaf_96_clk _00454_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[414\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06515__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ clknet_leaf_70_clk _00385_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[345\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11487__SET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07166__S0 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08283__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05489__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11425_ clknet_leaf_85_clk _00937_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07243__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09783__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ clknet_leaf_41_clk _00868_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[828\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11495__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08820__C net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ _02485_ net1493 net236 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
X_11287_ clknet_leaf_21_clk _00799_ net1182 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[759\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05518__A _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ net1126 net1454 net911 _05227_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__a31o_1
XANTENNA__06349__A2 _02451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1030 net1033 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_37_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_2
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10169_ net127 net917 net906 net1517 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a22o_1
XANTENNA__11101__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1063 net1064 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1074 core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_4
XANTENNA__07292__X _03397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09424__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1085 net1090 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_4
XFILLER_0_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1096 net1103 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06506__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05253__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_44_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06400_ net946 core.register_file.registers_state\[193\] net704 core.register_file.registers_state\[225\]
+ net643 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ net977 _03483_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06331_ net1032 _02431_ _02435_ net1006 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06904__S0 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09050_ net2167 net429 _05006_ net1002 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__a22o_1
X_06262_ core.register_file.registers_state\[4\] net710 net646 _02366_ vssd1 vssd1
+ vccd1 vccd1 _02367_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_59_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08001_ _03893_ _04085_ _04087_ _04079_ net492 net477 vssd1 vssd1 vccd1 vccd1 _04106_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10712__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06193_ net940 core.register_file.registers_state\[838\] net1013 vssd1 vssd1 vccd1
+ vccd1 _02298_ sky130_fd_sc_hd__a21o_1
XANTENNA__10369__A0 _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11838__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_102_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold502 core.register_file.registers_state\[682\] vssd1 vssd1 vccd1 vccd1 net1821
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold513 core.register_file.registers_state\[650\] vssd1 vssd1 vccd1 vccd1 net1832
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 core.register_file.registers_state\[233\] vssd1 vssd1 vccd1 vccd1 net1843
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06037__B2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09774__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold535 core.register_file.registers_state\[687\] vssd1 vssd1 vccd1 vccd1 net1854
+ sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap254 _04683_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_1
Xhold546 core.register_file.registers_state\[426\] vssd1 vssd1 vccd1 vccd1 net1865
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold557 core.register_file.registers_state\[538\] vssd1 vssd1 vccd1 vccd1 net1876
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold568 core.register_file.registers_state\[424\] vssd1 vssd1 vccd1 vccd1 net1887
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ core.IO_mod.data_from_mem\[8\] core.CPU_DAT_O\[8\] net801 vssd1 vssd1 vccd1
+ vccd1 _01104_ sky130_fd_sc_hd__mux2_1
Xhold579 core.register_file.registers_state\[294\] vssd1 vssd1 vccd1 vccd1 net1898
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08903_ net569 _04908_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__and2_1
XANTENNA__09526__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06023__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ net1118 _05069_ net376 net1878 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__a22o_1
XANTENNA__07537__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 core.register_file.registers_state\[644\] vssd1 vssd1 vccd1 vccd1 net2521
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ core.IO_mod.data_from_mem\[31\] core.IO_mod.input_reg\[31\] net250 vssd1
+ vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__mux2_1
XANTENNA__06958__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1213 core.register_file.registers_state\[855\] vssd1 vssd1 vccd1 vccd1 net2532
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A _01368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 core.register_file.registers_state\[728\] vssd1 vssd1 vccd1 vccd1 net2543
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 core.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05643__S0 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ net733 _04287_ _04756_ _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__o211a_4
XANTENNA__11218__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05977_ net1025 _02078_ _02081_ net717 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout462_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08458__B net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__RESET_B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ net498 _03670_ _03663_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_101_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08498__C1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ core.IO_mod.data_from_mem\[9\] net246 _04761_ vssd1 vssd1 vccd1 vccd1 _04762_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07647_ net506 _03703_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout727_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07170__C1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07578_ _01626_ _03620_ _03616_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__o21ai_4
XANTENNA__05720__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07148__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ _04943_ net420 net333 net2212 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06529_ _02630_ _02632_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1257_X net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10072__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ core.register_file.registers_state\[315\] net474 net544 vssd1 vssd1 vccd1
+ vccd1 _05040_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08761__X _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09214__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _04963_ net357 net425 net1714 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08921__B net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11210_ clknet_leaf_106_clk _00722_ net1139 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[682\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06281__X _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09765__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06123__S1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07096__Y _03201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11141_ clknet_leaf_87_clk _00653_ net1229 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[613\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06984__C1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XANTENNA__09517__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ clknet_leaf_60_clk _00584_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[544\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_37_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__07528__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ net724 _01778_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__and2_2
XANTENNA__07553__A _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05634__S0 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06169__A core.decoder.inst\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10565__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10925_ clknet_leaf_2_clk _00437_ net1139 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[397\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07700__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06456__X _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ clknet_leaf_13_clk _00368_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[328\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05711__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10735__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09453__A1 _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ clknet_leaf_66_clk _00299_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[259\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07464__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08671__X _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09205__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08831__B _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output91_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09419__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ clknet_leaf_105_clk _00920_ net1157 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[880\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09756__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06191__X _02296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__RESET_B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08964__B1 _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11339_ clknet_leaf_108_clk _00851_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[811\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07447__B net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__A _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06351__B _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__B1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05900_ net951 core.register_file.registers_state\[975\] net709 core.register_file.registers_state\[1007\]
+ net929 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06880_ net991 core.register_file.registers_state\[78\] net877 core.register_file.registers_state\[110\]
+ net824 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a221o_1
XANTENNA__06727__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07463__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05831_ net627 _01934_ _01935_ net717 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a31o_1
XANTENNA__08731__A3 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ core.pc.current_pc\[28\] _04603_ core.pc.current_pc\[29\] vssd1 vssd1 vccd1
+ vccd1 _04628_ sky130_fd_sc_hd__a21oi_1
X_05762_ _01408_ _01409_ core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o21a_4
XANTENNA__09141__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07501_ net772 _03594_ _03605_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__a21boi_1
X_08481_ _01710_ _04564_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__nand2_1
X_05693_ net629 _01794_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__or3_1
XFILLER_0_134_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07432_ _02534_ _02598_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06050__S0 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ core.register_file.registers_state\[538\] core.register_file.registers_state\[570\]
+ net868 vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11470__SET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09102_ net2237 net363 net351 _04845_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__a22o_1
X_06314_ net964 _02413_ _02418_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a21oi_1
X_07294_ _03142_ _03398_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__and2_1
XANTENNA__06018__S net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10048__B net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06245_ net1059 core.register_file.registers_state\[740\] net754 _02349_ vssd1 vssd1
+ vccd1 vccd1 _02350_ sky130_fd_sc_hd__a31o_1
X_09033_ net614 net217 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout210_A _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A _05063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold310 core.register_file.registers_state\[912\] vssd1 vssd1 vccd1 vccd1 net1629
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09747__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06176_ core.register_file.registers_state\[6\] net698 net640 _02280_ vssd1 vssd1
+ vccd1 vccd1 _02281_ sky130_fd_sc_hd__o211a_1
Xhold321 core.register_file.registers_state\[266\] vssd1 vssd1 vccd1 vccd1 net1640
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 net107 vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 core.register_file.registers_state\[274\] vssd1 vssd1 vccd1 vccd1 net1662
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 core.register_file.registers_state\[278\] vssd1 vssd1 vccd1 vccd1 net1673
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 core.register_file.registers_state\[881\] vssd1 vssd1 vccd1 vccd1 net1684
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold376 core.register_file.registers_state\[619\] vssd1 vssd1 vccd1 vccd1 net1695
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1217_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 core.register_file.registers_state\[285\] vssd1 vssd1 vccd1 vccd1 net1706
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _05090_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_2
XANTENNA__06430__A1 core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold398 core.register_file.registers_state\[304\] vssd1 vssd1 vccd1 vccd1 net1717
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ core.decoder.inst\[24\] core.CPU_DAT_O\[24\] net891 vssd1 vssd1 vccd1 vccd1
+ _01088_ sky130_fd_sc_hd__mux2_1
Xfanout812 net815 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_4
Xfanout823 _01459_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_4
Xfanout834 net838 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08707__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 net861 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
X_09866_ _04939_ net388 net268 net1871 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__a22o_1
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1005_X net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10608__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout878 net882 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_2
Xhold1010 core.register_file.registers_state\[54\] vssd1 vssd1 vccd1 vccd1 net2329
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1021 core.register_file.registers_state\[112\] vssd1 vssd1 vccd1 vccd1 net2340
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07373__A _03475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05445__X _01550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout889 net890 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__buf_4
XANTENNA__09380__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ core.IO_mod.data_from_mem\[28\] net246 _04863_ vssd1 vssd1 vccd1 vccd1 _04864_
+ sky130_fd_sc_hd__a21o_1
Xhold1032 core.register_file.registers_state\[752\] vssd1 vssd1 vccd1 vccd1 net2351
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 core.register_file.registers_state\[755\] vssd1 vssd1 vccd1 vccd1 net2362
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1054 core.register_file.registers_state\[763\] vssd1 vssd1 vccd1 vccd1 net2373
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _04807_ net387 net271 net1835 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 core.register_file.registers_state\[711\] vssd1 vssd1 vccd1 vccd1 net2384
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 core.register_file.registers_state\[576\] vssd1 vssd1 vccd1 vccd1 net2395
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 core.register_file.registers_state\[80\] vssd1 vssd1 vccd1 vccd1 net2406
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ net608 net217 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 core.register_file.registers_state\[498\] vssd1 vssd1 vccd1 vccd1 net2417
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09132__A0 _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ net568 net607 _04746_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06497__A1 _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ clknet_leaf_59_clk _00222_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[182\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07694__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10293__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06276__X _02381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ clknet_leaf_76_clk net1513 net1260 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ clknet_leaf_72_clk _00153_ net1272 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10572_ clknet_leaf_102_clk _00084_ net1162 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08932__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09199__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09738__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05994__C net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ clknet_leaf_57_clk _00636_ net1297 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[596\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11055_ clknet_leaf_83_clk _00567_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[527\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05355__X _01460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07283__A _03289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09371__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ net1587 net540 net519 _05103_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__a22o_1
XANTENNA__06185__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07921__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07921__B2 _03972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05932__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09123__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09702__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08477__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07134__C1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__B _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06032__S0 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ clknet_leaf_42_clk _00420_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06488__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11888_ clknet_leaf_50_clk _01357_ net1307 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06627__A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09003__A _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09426__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839_ clknet_leaf_20_clk _00351_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[311\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09497__X _05060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07988__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06030_ net620 _02133_ _02134_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__and3_1
XANTENNA__06660__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09729__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06412__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ net504 _03645_ _03783_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09720_ _04912_ net293 net277 net2290 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__a22o_1
X_06932_ net986 core.register_file.registers_state\[459\] net862 core.register_file.registers_state\[491\]
+ net978 vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09362__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _04737_ net294 net285 net1755 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__a22o_1
X_06863_ _02966_ _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06176__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ _04186_ _04200_ _04215_ _04255_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__or4_1
XANTENNA__06271__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05814_ core.register_file.registers_state\[274\] core.register_file.registers_state\[306\]
+ core.register_file.registers_state\[402\] core.register_file.registers_state\[434\]
+ net714 net1021 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__mux4_1
X_09582_ _04929_ net400 net300 net1814 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06794_ net968 _02895_ _02898_ _02889_ _02892_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09114__A0 _04730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08533_ _01385_ net553 net574 vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__mux2_1
X_05745_ net1063 core.register_file.registers_state\[84\] core.register_file.registers_state\[116\]
+ net691 net649 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07125__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__B net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout258_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08464_ _04548_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__xnor2_1
X_05676_ net554 _01778_ _01779_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07415_ core.register_file.registers_state\[984\] core.register_file.registers_state\[1016\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09417__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__A _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08395_ _04485_ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout425_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1167_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07428__B1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07346_ _03449_ _03450_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11275__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06326__S1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05439__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11406__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06100__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ net769 _03374_ _03381_ _03368_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a31o_4
XFILLER_0_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08640__A2 _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ net742 net462 _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__and3_1
XANTENNA__07368__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06228_ core.register_file.registers_state\[517\] net698 net639 _02332_ vssd1 vssd1
+ vccd1 vccd1 _02333_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout794_A _01455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold140 core.register_file.registers_state\[29\] vssd1 vssd1 vccd1 vccd1 net1459
+ sky130_fd_sc_hd__dlygate4sd3_1
X_06159_ _02260_ _02261_ _02262_ _02263_ net929 net964 vssd1 vssd1 vccd1 vccd1 _02264_
+ sky130_fd_sc_hd__mux4_1
Xhold151 core.register_file.registers_state\[12\] vssd1 vssd1 vccd1 vccd1 net1470
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_X net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold162 core.CPU_DAT_I\[31\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 net142 vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold184 net118 vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08306__A1_N _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 net177 vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05319__C core.decoder.inst\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout961_A _01373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout620 net621 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout631 net632 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09918_ core.decoder.inst\[7\] core.CPU_DAT_O\[7\] net892 vssd1 vssd1 vccd1 vccd1
+ _01071_ sky130_fd_sc_hd__mux2_1
Xfanout642 _01516_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_8
Xfanout653 net664 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 _01515_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout675 net676 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09353__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout686 net687 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout697 net701 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_4
X_09849_ _04905_ net389 net267 net1863 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__a22o_1
XANTENNA__10241__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__C1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08927__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ clknet_leaf_76_clk _01312_ net1261 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10153__B1_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08646__B net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07667__A0 _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ clknet_leaf_36_clk _01254_ net1221 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07550__B _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05351__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ clknet_leaf_36_clk _01185_ net1221 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09408__A1 _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ clknet_leaf_52_clk _00136_ net1303 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07419__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11086__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__X _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10555_ clknet_leaf_25_clk _00067_ net1186 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07278__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net1422 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10998__RESET_B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09592__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ clknet_leaf_67_clk _00619_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[579\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09344__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11038_ clknet_leaf_97_clk _00550_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[510\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09895__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08837__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09647__A1 _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05381__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__C1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05530_ core.register_file.registers_state\[26\] core.register_file.registers_state\[58\]
+ core.register_file.registers_state\[154\] core.register_file.registers_state\[186\]
+ net696 net653 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05669__C1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05261__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05461_ _01562_ _01564_ _01565_ net933 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06330__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07200_ _03302_ _03304_ net770 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__a21o_1
XANTENNA__06881__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ _03686_ _04244_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__o21ba_2
X_05392_ core.decoder.inst\[14\] _01417_ _01425_ _01489_ vssd1 vssd1 vccd1 vccd1 _01497_
+ sky130_fd_sc_hd__or4b_1
XANTENNA__06791__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06308__S1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07131_ _03235_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__inv_2
XANTENNA__08083__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11579__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07188__A _03289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07062_ net1107 core.register_file.registers_state\[679\] core.register_file.registers_state\[647\]
+ net848 net808 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__a221o_1
XANTENNA__06092__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput201 net201 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_3_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06013_ core.register_file.registers_state\[555\] core.register_file.registers_state\[523\]
+ net668 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
XANTENNA__05841__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08386__B2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09583__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06397__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07964_ _01365_ _02084_ _02931_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05436__A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09335__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ net205 core.register_file.registers_state\[727\] net278 vssd1 vssd1 vccd1
+ vccd1 _00767_ sky130_fd_sc_hd__mux2_1
X_06915_ _03018_ _03019_ net1086 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__o21a_1
XANTENNA__10061__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07895_ net579 _03998_ _03999_ _03995_ _03997_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__a311o_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _05007_ net396 net391 net2166 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__a22o_1
X_06846_ core.register_file.registers_state\[687\] core.register_file.registers_state\[655\]
+ net853 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05870__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ net241 net2085 net305 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout542_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06777_ core.register_file.registers_state\[272\] core.register_file.registers_state\[304\]
+ core.register_file.registers_state\[400\] core.register_file.registers_state\[432\]
+ net865 net1073 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1284_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ _01633_ _04595_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05728_ core.register_file.registers_state\[788\] core.register_file.registers_state\[820\]
+ core.register_file.registers_state\[916\] core.register_file.registers_state\[948\]
+ net713 net1023 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__mux4_1
XANTENNA__11456__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ _05020_ net320 net262 net1676 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08447_ _04515_ _04533_ _04524_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05602__C _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05659_ _01762_ _01763_ net719 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1072_X net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A _01460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06872__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__A _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ _02017_ _04469_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05321__D net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08074__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ net1095 core.register_file.registers_state\[731\] core.register_file.registers_state\[763\]
+ net836 net818 vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09810__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10340_ _02485_ net1464 net233 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10946__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10271_ net2 net903 net795 net2529 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_72_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09574__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06730__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout450 _02530_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_2
XANTENNA__08129__B2 _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout461 _05060_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_4
Xfanout472 _05127_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 _02516_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09877__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout494 net496 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07337__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06235__S0 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07561__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05899__C1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11725_ clknet_leaf_47_clk _01237_ net1306 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08663__Y _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ clknet_leaf_47_clk _01168_ net1306 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11721__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ clknet_leaf_82_clk _00119_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_11587_ clknet_leaf_26_clk _01099_ net1203 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09801__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09000__B _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07812__B1 _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ clknet_leaf_107_clk _00050_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold909 core.register_file.registers_state\[247\] vssd1 vssd1 vccd1 vccd1 net2228
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10469_ net1338 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09565__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09427__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10175__B2 core.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09317__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05256__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ net1097 core.register_file.registers_state\[339\] core.register_file.registers_state\[371\]
+ net840 net980 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07680_ net449 net550 net441 net501 vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__o31a_1
XANTENNA__08540__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06777__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06631_ net1105 core.register_file.registers_state\[85\] core.register_file.registers_state\[117\]
+ net851 net811 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__o221a_1
XANTENNA__11251__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05354__B2 _01395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09350_ net1119 _04998_ net415 net1718 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10819__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06562_ core.register_file.registers_state\[535\] core.register_file.registers_state\[567\]
+ net868 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XANTENNA__09096__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08301_ _04386_ _04390_ _04399_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05513_ _01493_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__nor2_1
X_09281_ net2187 _04891_ net337 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
X_06493_ net555 _02597_ _02563_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07500__C1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08232_ _01380_ net577 vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__nor2_1
X_05444_ _01527_ _01534_ _01542_ _01548_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__o22a_4
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07410__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ _04260_ _04261_ _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10337__A _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05375_ net975 _01478_ _01479_ net1068 _01477_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__o311a_1
XFILLER_0_126_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10849__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07114_ core.register_file.registers_state\[37\] net842 vssd1 vssd1 vccd1 vccd1 _03219_
+ sky130_fd_sc_hd__or2_1
X_08094_ _03831_ _04063_ net534 vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10056__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload60 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_110_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07045_ core.register_file.registers_state\[7\] net878 net808 _03149_ vssd1 vssd1
+ vccd1 vccd1 _03150_ sky130_fd_sc_hd__o211a_1
Xclkload71 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__09845__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload82 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout1032_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09556__A0 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__07646__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09020__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__B2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ net2420 net429 _04970_ net1000 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09308__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ net1003 _04050_ _04051_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07319__C1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05593__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07878_ net507 _03675_ _03652_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__o21ai_1
XANTENNA__05316__D net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09617_ _04988_ net395 net391 net1615 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__a22o_1
X_06829_ _02084_ _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_104_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout924_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1287_X net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ net221 net2248 net304 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__mux2_1
XANTENNA__08764__X _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09087__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09479_ _04989_ net323 net263 net1830 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08924__B net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11510_ clknet_leaf_61_clk _01022_ net1281 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[982\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06845__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ clknet_leaf_81_clk _00953_ net1255 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[913\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09795__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ clknet_leaf_103_clk _00884_ net1156 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[844\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08062__A3 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10323_ _05108_ net1580 net238 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input53_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ net1125 net1463 net910 _05235_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__a31o_1
XANTENNA__08004__X _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09011__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1213 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__buf_2
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10185_ net113 net917 net907 net1572 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a22o_1
XANTENNA__08939__X _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06230__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1245 net1246 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_2
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1267 net1268 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_2
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_8
Xfanout1278 net1314 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout291 _05080_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
Xfanout1289 net1292 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11378__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05363__X _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__RESET_B net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09078__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09710__S net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07628__A3 _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ clknet_leaf_76_clk net1730 net1261 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11639_ clknet_leaf_72_clk _01151_ net1269 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10157__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08589__A1 core.decoder.inst\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09786__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08850__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold706 core.register_file.registers_state\[517\] vssd1 vssd1 vccd1 vccd1 net2025
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold717 core.register_file.registers_state\[512\] vssd1 vssd1 vccd1 vccd1 net2036
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07261__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold728 core.register_file.registers_state\[255\] vssd1 vssd1 vccd1 vccd1 net2047
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold739 core.register_file.registers_state\[312\] vssd1 vssd1 vccd1 vccd1 net2058
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09538__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09002__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11617__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07013__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05257__Y _01372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ net741 _04751_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07013__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ _03749_ _03754_ net485 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06221__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08781_ net570 net610 net213 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__and3_1
X_05993_ net1049 core.register_file.registers_state\[172\] net675 core.register_file.registers_state\[140\]
+ net640 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a221o_1
X_07732_ _03657_ _03834_ _03836_ _03832_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07913__B _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__A2 _03412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09710__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05714__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _03715_ _03725_ net506 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux2_1
X_09402_ net2476 net224 net407 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__mux2_1
X_06614_ _01781_ _02687_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__xnor2_1
X_07594_ net453 _03052_ net445 net502 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ net1119 net464 _04964_ net414 net1690 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06545_ net975 _02648_ _02649_ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout338_A _05046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06288__C1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05720__Y _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09264_ net2249 net223 net338 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06476_ _02579_ _02580_ net958 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06545__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08215_ _04004_ _04043_ _04298_ _04319_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__or4b_1
XFILLER_0_118_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05427_ core.register_file.registers_state\[926\] core.register_file.registers_state\[958\]
+ net700 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09195_ _04995_ net359 net425 net1728 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout505_A _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1247_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09777__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ net488 _04133_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__nand2_1
X_05358_ net1067 _01397_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__nand2_4
XFILLER_0_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08760__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ net500 _03722_ _03727_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a21bo_1
X_05289_ core.control_logic.instruction\[5\] core.control_logic.instruction\[6\] vssd1
+ vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07028_ core.register_file.registers_state\[776\] core.register_file.registers_state\[808\]
+ core.register_file.registers_state\[904\] core.register_file.registers_state\[936\]
+ net874 net1070 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_8_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout874_A _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07004__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__B1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1202_X net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08759__X _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06212__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 core.register_file.registers_state\[931\] vssd1 vssd1 vccd1 vccd1 net1330
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 core.register_file.registers_state\[943\] vssd1 vssd1 vccd1 vccd1 net1341
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 core.register_file.registers_state\[946\] vssd1 vssd1 vccd1 vccd1 net1352
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold44 core.register_file.registers_state\[930\] vssd1 vssd1 vccd1 vccd1 net1363
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ net2296 net368 _04959_ net433 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 core.register_file.registers_state\[944\] vssd1 vssd1 vccd1 vccd1 net1374
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 core.register_file.registers_state\[965\] vssd1 vssd1 vccd1 vccd1 net1385
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07823__B _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 core.register_file.registers_state\[990\] vssd1 vssd1 vccd1 vccd1 net1396
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06279__X _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold88 core.register_file.registers_state\[948\] vssd1 vssd1 vccd1 vccd1 net1407
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 core.register_file.registers_state\[16\] vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08504__A1 _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__A0 _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ clknet_leaf_19_clk _00453_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[413\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11400__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10872_ clknet_leaf_5_clk _00384_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[344\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08935__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10075__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07166__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09480__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07491__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07491__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11424_ clknet_leaf_56_clk _00936_ net1294 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09232__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11355_ clknet_leaf_21_clk _00867_ net1190 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07286__A _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _02514_ net1458 net236 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
XANTENNA__06451__C1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11286_ clknet_leaf_59_clk _00798_ net1287 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[758\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ net80 net921 vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10664__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09940__A0 core.decoder.inst\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1020 net1024 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_4
Xfanout1031 net1032 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_4
XANTENNA__09705__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1042 net1053 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__buf_2
Xfanout1053 core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_4
X_10168_ net126 net916 net907 net1659 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a22o_1
XANTENNA__05557__A1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06754__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__buf_2
XANTENNA__08829__B _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_4
Xfanout1086 net1087 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
Xfanout1097 net1099 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_10099_ _04317_ net557 net588 core.pc.current_pc\[19\] net471 vssd1 vssd1 vccd1 vccd1
+ _05159_ sky130_fd_sc_hd__o221a_1
XANTENNA__09299__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09006__A _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08259__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_108_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10066__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06330_ _02432_ _02433_ net965 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06809__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06809__B2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09471__A2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06261_ net952 core.register_file.registers_state\[36\] net765 vssd1 vssd1 vccd1
+ vccd1 _02366_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08000_ _04079_ _04085_ net484 vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__mux2_1
XANTENNA__09759__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06690__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08580__A core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06192_ core.register_file.registers_state\[806\] core.register_file.registers_state\[774\]
+ core.register_file.registers_state\[934\] core.register_file.registers_state\[902\]
+ net675 net1014 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__mux4_1
XANTENNA__09223__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07234__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 core.register_file.registers_state\[427\] vssd1 vssd1 vccd1 vccd1 net1822
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 core.register_file.registers_state\[883\] vssd1 vssd1 vccd1 vccd1 net1833
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold525 core.register_file.registers_state\[393\] vssd1 vssd1 vccd1 vccd1 net1844
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap244 _04703_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
Xhold536 core.register_file.registers_state\[909\] vssd1 vssd1 vccd1 vccd1 net1855
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold547 core.register_file.registers_state\[514\] vssd1 vssd1 vccd1 vccd1 net1866
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09951_ net1574 core.CPU_DAT_O\[7\] net798 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
Xhold558 core.register_file.registers_state\[575\] vssd1 vssd1 vccd1 vccd1 net1877
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05709__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold569 core.register_file.registers_state\[783\] vssd1 vssd1 vccd1 vccd1 net1888
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06993__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ _04741_ net602 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ net1118 _05068_ net376 net1862 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__a22o_1
XANTENNA__07537__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09931__A0 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ net2366 net468 net436 _04877_ vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__a22o_1
Xhold1203 core.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05548__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1214 core.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11229__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1225 core.register_file.registers_state\[203\] vssd1 vssd1 vccd1 vccd1 net2544
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout288_A _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1236 core.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ core.IO_mod.data_from_mem\[20\] net247 _04818_ vssd1 vssd1 vccd1 vccd1 _04819_
+ sky130_fd_sc_hd__a21o_2
XANTENNA__05643__S1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06099__X _02204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05976_ net1004 _02079_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__or3_1
X_07715_ net510 _03819_ _03818_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__a21oi_1
X_08695_ core.IO_mod.input_reg\[9\] net250 net725 vssd1 vssd1 vccd1 vccd1 _04761_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_101_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout455_A _02529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07646_ net491 _03750_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08755__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07577_ net1003 _03612_ net580 _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout622_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_X net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10057__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07148__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ _04941_ net420 net333 net2326 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a22o_1
XANTENNA__09998__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06528_ _02630_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__nor2_1
XANTENNA__09462__A2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ net558 _04857_ _05039_ net339 net1999 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06459_ net1035 net747 core.register_file.registers_state\[792\] vssd1 vssd1 vccd1
+ vccd1 _02564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05610__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07658__X _03763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ _04704_ net1958 net426 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__mux2_1
XANTENNA__09214__A2 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout991_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08921__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _03383_ _04231_ _04233_ _03382_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__o22a_1
XANTENNA__07225__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10687__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11140_ clknet_leaf_81_clk _00652_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[612\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08973__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11071_ clknet_leaf_15_clk _00583_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[543\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XANTENNA__07528__A2 _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__A0 core.decoder.inst\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ net1495 net542 net521 _05111_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_78_clk_X clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05539__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05539__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__B _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06200__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05634__S1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06169__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ clknet_leaf_102_clk _00436_ net1162 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09260__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07700__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10855_ clknet_leaf_93_clk _00367_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[327\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_16_clk_X clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10786_ clknet_leaf_78_clk _00298_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[258\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09453__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05475__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09205__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07216__A1 _01506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ clknet_leaf_79_clk _00919_ net1253 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[879\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08413__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05529__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11338_ clknet_leaf_107_clk _00850_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[810\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08964__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05778__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05778__B2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ clknet_leaf_87_clk _00781_ net1229 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[741\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07744__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08192__A2 _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05830_ net654 _01933_ _01932_ net616 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_59_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05264__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05761_ _01825_ _01826_ _01862_ _01863_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
X_07500_ net780 _03599_ _03604_ net768 vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__o211ai_1
X_08480_ _01383_ net552 net574 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__mux2_1
X_05692_ _01786_ _01796_ _01795_ net1019 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_134_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07431_ net771 _03523_ _03534_ _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a22o_4
XANTENNA__06050__S1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07362_ net1082 _03463_ _03466_ net1066 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09444__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09101_ net2535 net363 net352 _04839_ vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__a22o_1
X_06313_ net1031 _02415_ _02417_ net934 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07293_ _03139_ _03141_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__or2_1
XANTENNA__08581__Y _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05466__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09032_ net1907 net427 _04994_ net998 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__a22o_1
XANTENNA__07919__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06663__C1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06244_ net952 core.register_file.registers_state\[708\] vssd1 vssd1 vccd1 vccd1
+ _02349_ sky130_fd_sc_hd__and2_1
XANTENNA__08514__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06382__X _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07207__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold300 _01114_ vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold311 core.register_file.registers_state\[399\] vssd1 vssd1 vccd1 vccd1 net1630
+ sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ net941 core.register_file.registers_state\[38\] net761 vssd1 vssd1 vccd1
+ vccd1 _02280_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold322 core.register_file.registers_state\[283\] vssd1 vssd1 vccd1 vccd1 net1641
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06415__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold333 core.register_file.registers_state\[397\] vssd1 vssd1 vccd1 vccd1 net1652
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 core.register_file.registers_state\[391\] vssd1 vssd1 vccd1 vccd1 net1663
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 core.register_file.registers_state\[814\] vssd1 vssd1 vccd1 vccd1 net1674
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold366 core.register_file.registers_state\[546\] vssd1 vssd1 vccd1 vccd1 net1685
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10064__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06261__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 core.register_file.registers_state\[914\] vssd1 vssd1 vccd1 vccd1 net1696
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold388 core.register_file.registers_state\[300\] vssd1 vssd1 vccd1 vccd1 net1707
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net804 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
X_09934_ net1005 core.CPU_DAT_O\[23\] net893 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XANTENNA__06430__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold399 core.register_file.registers_state\[402\] vssd1 vssd1 vccd1 vccd1 net1718
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1112_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 net815 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout824 net826 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_4
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 _01458_ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_4
XANTENNA__09904__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ net559 _04937_ net458 net269 net1833 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__a32o_1
Xfanout857 net861 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__buf_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 core.register_file.registers_state\[688\] vssd1 vssd1 vccd1 vccd1 net2319
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net874 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
XANTENNA_fanout572_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1011 core.register_file.registers_state\[864\] vssd1 vssd1 vccd1 vccd1 net2330
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 net882 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_4
Xhold1022 core.register_file.registers_state\[467\] vssd1 vssd1 vccd1 vccd1 net2341
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ core.IO_mod.input_reg\[28\] net250 net726 vssd1 vssd1 vccd1 vccd1 _04863_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09380__B2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06813__S0 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1033 core.register_file.registers_state\[668\] vssd1 vssd1 vccd1 vccd1 net2352
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 core.register_file.registers_state\[861\] vssd1 vssd1 vccd1 vccd1 net2363
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _04802_ net385 net273 net1808 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__a22o_1
XANTENNA__11335__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1055 core.register_file.registers_state\[602\] vssd1 vssd1 vccd1 vccd1 net2374
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 core.register_file.registers_state\[190\] vssd1 vssd1 vccd1 vccd1 net2385
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net733 _04043_ net526 _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__o211a_4
XANTENNA_clkbuf_leaf_90_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 core.register_file.registers_state\[310\] vssd1 vssd1 vccd1 vccd1 net2396
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1088 core.register_file.registers_state\[164\] vssd1 vssd1 vccd1 vccd1 net2407
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05959_ _02062_ _02063_ net1025 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1099 core.register_file.registers_state\[344\] vssd1 vssd1 vccd1 vccd1 net2418
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout837_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10278__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ net606 _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__and2_1
XANTENNA__07143__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07629_ _03615_ _03626_ _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06497__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11485__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ clknet_leaf_107_clk _00152_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08772__X _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09435__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__B net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10571_ clknet_leaf_109_clk _00083_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08932__B net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05457__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06406__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08946__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ clknet_leaf_11_clk _00635_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[595\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ clknet_leaf_82_clk _00566_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[526\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10005_ net724 _02083_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_30_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06185__A1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07921__A2 _04016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07851__X _03956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__C_N _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05932__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_101_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05812__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07685__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08882__A0 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ clknet_leaf_25_clk _00419_ net1185 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[379\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06032__S1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11887_ clknet_leaf_50_clk _01356_ net1308 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09778__X _05085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09003__B _04751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10838_ clknet_leaf_59_clk _00350_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08682__X _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10769_ clknet_leaf_73_clk _00281_ net1272 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[241\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05259__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06948__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06412__A2 _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07980_ _03640_ _03641_ net508 vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__mux2_1
XANTENNA__11358__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06931_ net986 core.register_file.registers_state\[331\] net862 core.register_file.registers_state\[363\]
+ net1069 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a221o_1
XANTENNA__09362__A1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09650_ _04731_ net294 net285 net2434 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__a22o_1
X_06862_ _02962_ _02965_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__nor2_1
X_08601_ _03839_ _04672_ _04675_ _03862_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__or4b_1
XANTENNA__07761__X _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05813_ _01914_ _01917_ net635 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a21oi_1
X_09581_ _04927_ net400 net300 net2343 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__a22o_1
X_06793_ net805 _02896_ _02897_ net1084 vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a211o_1
XANTENNA__06271__S1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05923__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ core.pc.current_pc\[27\] _04611_ net595 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05744_ _01846_ _01848_ net623 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a21o_1
XANTENNA__08509__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09665__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07413__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05722__A _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _04531_ _04535_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__nor2_1
XANTENNA__08873__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05675_ net585 _01764_ _01777_ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ core.register_file.registers_state\[856\] core.register_file.registers_state\[888\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__mux2_1
XANTENNA__06884__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08394_ _04470_ _04475_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10059__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07345_ _03446_ _03448_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1062_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _05029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06636__C1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06100__A1 core.decoder.inst\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ net787 _03377_ _03380_ net782 vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__a211o_1
XANTENNA__08640__A3 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ net612 _04775_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06227_ core.register_file.registers_state\[549\] net675 vssd1 vssd1 vccd1 vccd1
+ _02332_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 core.register_file.registers_state\[961\] vssd1 vssd1 vccd1 vccd1 net1449
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 core.IO_mod.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ core.register_file.registers_state\[807\] core.register_file.registers_state\[775\]
+ net682 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
Xhold152 core.IO_mod.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06939__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold163 _01232_ vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold174 net193 vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _01226_ vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
X_06089_ core.register_file.registers_state\[73\] core.register_file.registers_state\[105\]
+ net699 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XANTENNA__05319__D net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1115_X net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 net146 vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _04669_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
Xfanout621 net626 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09917_ core.control_logic.instruction\[6\] core.CPU_DAT_O\[6\] net891 vssd1 vssd1
+ vccd1 vccd1 _01070_ sky130_fd_sc_hd__mux2_1
Xfanout632 _01521_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_70_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout643 net645 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_4
Xfanout654 net656 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_4
XANTENNA_fanout954_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout665 net666 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_97_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout676 net679 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _04903_ net389 net267 net1916 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__a22o_1
Xfanout687 net689 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout698 net701 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06167__B2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__X _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08561__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ net1121 net605 net383 vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_83_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ clknet_leaf_52_clk _01311_ net1303 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07116__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09656__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05632__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ clknet_leaf_36_clk _01253_ net1221 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07667__A1 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11672_ clknet_leaf_36_clk _01184_ net1221 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07419__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10623_ clknet_leaf_94_clk _00135_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ clknet_leaf_8_clk _00066_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07278__B _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10485_ net1415 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05850__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08919__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09041__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A1 _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ clknet_leaf_80_clk _00618_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[578\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05807__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09344__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ clknet_leaf_18_clk _00549_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[509\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08677__X _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__B1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05366__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08837__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09647__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06638__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05542__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__A0 _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05460_ core.register_file.registers_state\[797\] core.register_file.registers_state\[829\]
+ core.register_file.registers_state\[925\] core.register_file.registers_state\[957\]
+ net696 net1011 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05391_ core.control_logic.instruction\[4\] _01402_ _01404_ vssd1 vssd1 vccd1 vccd1
+ _01496_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
X_07130_ _03231_ _03233_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08064__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07061_ core.register_file.registers_state\[551\] core.register_file.registers_state\[519\]
+ net848 vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__mux2_1
XANTENNA__07830__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11180__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput202 net202 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__07756__X _03861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06012_ _02115_ _02116_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07043__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10193__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07408__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _02084_ _02931_ net578 vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_79_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09335__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06914_ net1098 core.register_file.registers_state\[460\] core.register_file.registers_state\[492\]
+ net841 net1075 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__o221a_1
X_09702_ net213 net2019 net280 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07894_ _01827_ _02747_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__nand2_1
XANTENNA__09886__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07897__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06845_ net777 _02942_ _02949_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_65_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09633_ net2278 net393 _05077_ net1002 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout270_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout368_A _04898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09564_ net243 net2411 net305 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__mux2_1
X_06776_ net789 _02877_ _02880_ net775 vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__o211a_1
XANTENNA__09099__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ _01633_ _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__nor2_1
X_05727_ net930 _01830_ _01831_ net965 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a31o_1
XANTENNA__10248__A3 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _05018_ net326 net264 net1720 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1277_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ _01896_ _04511_ _04525_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05658_ net1030 _01748_ _01749_ _01752_ net1006 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06321__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06321__B2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08377_ _02017_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_119_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05589_ net1026 _01689_ _01692_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout702_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1065_X net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06609__C1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07328_ net780 _03430_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08074__A1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06283__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06085__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07259_ net1089 _03361_ _03363_ net1080 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1232_X net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07666__X _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ core.BUSY_O net905 wb.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_72_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11673__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10184__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__B1 _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout440 _04713_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_4
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 net455 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout462 net465 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_6
Xfanout473 _05127_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08938__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09877__A2 _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06235__S1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08657__B _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05899__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06458__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11724_ clknet_leaf_48_clk _01236_ net1306 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08673__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06312__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ clknet_leaf_47_clk _01167_ net1306 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10606_ clknet_leaf_89_clk _00118_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_11586_ clknet_leaf_26_clk _01098_ net1203 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07812__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__C1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10537_ clknet_leaf_39_clk _00049_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05823__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10468_ net1364 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06921__A _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07025__C1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ net1459 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06379__A1 _01375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06379__B2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10175__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09009__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05537__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05587__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09868__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06000__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ core.register_file.registers_state\[21\] core.register_file.registers_state\[53\]
+ net879 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06551__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06551__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06561_ net1082 _02665_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08300_ _04386_ _04390_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__or3_1
XANTENNA__08854__Y _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05512_ _01395_ _01403_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__or2_1
X_09280_ net2288 net214 net338 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
XANTENNA__06839__C1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06492_ _02581_ _02582_ _02590_ _02596_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__06303__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08583__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08231_ _01495_ _03740_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or2_4
X_05443_ _01546_ _01547_ net722 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _03657_ _03772_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05374_ net1100 core.register_file.registers_state\[862\] core.register_file.registers_state\[894\]
+ net843 net981 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__o221a_1
XANTENNA__09253__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06067__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07113_ net1098 core.register_file.registers_state\[133\] net841 core.register_file.registers_state\[165\]
+ net820 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o221a_1
X_08093_ net534 _04060_ _04197_ _03685_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_71_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload50 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_109_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07927__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ core.register_file.registers_state\[39\] net848 vssd1 vssd1 vccd1 vccd1 _03149_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload61 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_110_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06831__A _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload72 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_110_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload83 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload94 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_8
XFILLER_0_101_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10166__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05447__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ net743 net465 _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout485_A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ _02146_ _03052_ net578 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09859__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07877_ _03650_ _03798_ _03981_ _03730_ _03979_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__o221a_1
XANTENNA__08110__X _04215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09616_ net999 _04986_ net457 net392 net1647 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__a32o_1
X_06828_ _02114_ _02526_ net538 vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_104_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09547_ _04890_ net2320 net303 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__mux2_1
X_06759_ core.register_file.registers_state\[593\] core.register_file.registers_state\[625\]
+ net883 vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08295__A1 _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ _04987_ net315 net261 net1638 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__a22o_1
XANTENNA__05728__S0 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__RESET_B net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08924__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08429_ core.pc.current_pc\[18\] _04502_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05502__C1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08047__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11440_ clknet_leaf_104_clk _00952_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload0 clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_46_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09244__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10247__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06058__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ clknet_leaf_110_clk _00883_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[843\]
+ sky130_fd_sc_hd__dfrtp_1
X_10322_ _05107_ net1558 net237 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07837__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06741__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10253_ net88 net914 vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__and2_1
XANTENNA__07556__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05357__A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1202 net1209 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_2
XANTENNA_input46_A gpio_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ net1729 net916 net906 core.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 _01220_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11419__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1213 net1224 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_2
Xfanout1224 net1314 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1235 net1236 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 net1250 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__clkbuf_2
Xfanout1257 net1278 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06781__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1268 net1277 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 net273 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09263__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1279 net1281 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_4
Xfanout281 _05082_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_8
Xfanout292 net298 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05741__C1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09499__A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09483__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11347__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11707_ clknet_leaf_49_clk net1486 net1309 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11638_ clknet_leaf_49_clk _01150_ net1309 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09235__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08589__A2 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11569_ clknet_leaf_28_clk _01081_ net1194 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07797__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__B _04751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 core.register_file.registers_state\[764\] vssd1 vssd1 vccd1 vccd1 net2026
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold718 core.register_file.registers_state\[358\] vssd1 vssd1 vccd1 vccd1 net2037
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 core.register_file.registers_state\[776\] vssd1 vssd1 vccd1 vccd1 net2048
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10911__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11099__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ net265 _03898_ _03902_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06221__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07753__Y _03858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08780_ net610 net213 vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05992_ _02088_ _02089_ _02095_ _02096_ net960 net933 vssd1 vssd1 vccd1 vccd1 _02097_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08578__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07731_ net493 _03678_ _03835_ net513 vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07662_ net500 _03722_ _03766_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_133_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06524__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06613_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__inv_2
X_09401_ net2079 net225 net407 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__mux2_1
X_07593_ net453 _03080_ net445 net508 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a31o_1
XANTENNA__10936__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08584__Y _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__A1 core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06544_ net1104 core.register_file.registers_state\[860\] core.register_file.registers_state\[892\]
+ net850 net982 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__o221a_1
X_09332_ _04704_ net1982 net414 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__mux2_1
XANTENNA__09474__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10084__A1 _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06288__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ net2507 net224 net338 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06475_ net932 _02575_ _02576_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__or3_1
XANTENNA__07485__C1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_A _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08214_ _04028_ _04064_ _04259_ _04268_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05426_ net1048 core.register_file.registers_state\[990\] core.register_file.registers_state\[1022\]
+ net678 net1029 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__o221a_1
X_09194_ _04993_ net353 net423 net1623 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__a22o_1
XANTENNA__09226__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08145_ _02384_ _03260_ _03621_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__a31o_1
X_05357_ net968 net896 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__nor2_8
XFILLER_0_114_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout400_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05876__S net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08076_ net480 _04056_ _04118_ net491 vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__o211a_1
X_05288_ core.control_logic.instruction\[2\] core.control_logic.instruction\[3\] core.control_logic.instruction\[1\]
+ core.control_logic.instruction\[0\] vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__or4bb_2
XANTENNA__05799__C1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06561__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07027_ net971 _03130_ _03131_ _03129_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_8_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1028_X net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__X _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 core.register_file.registers_state\[932\] vssd1 vssd1 vccd1 vccd1 net1331
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06212__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 core.register_file.registers_state\[971\] vssd1 vssd1 vccd1 vccd1 net1342
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net567 net243 net736 vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__and3_1
Xhold34 core.register_file.registers_state\[958\] vssd1 vssd1 vccd1 vccd1 net1353
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 core.register_file.registers_state\[994\] vssd1 vssd1 vccd1 vccd1 net1364
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 core.register_file.registers_state\[945\] vssd1 vssd1 vccd1 vccd1 net1375
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 net138 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07929_ net579 _04032_ _04033_ _04031_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a31o_1
Xhold78 core.register_file.registers_state\[30\] vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05971__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 core.register_file.registers_state\[5\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10940_ clknet_leaf_40_clk _00452_ net1216 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[412\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06515__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06515__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ clknet_leaf_22_clk _00383_ net1181 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[343\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08935__B net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09465__A0 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10075__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09217__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08951__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07228__C1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11423_ clknet_leaf_62_clk _00935_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[895\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__B1 _03883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07567__A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ clknet_leaf_8_clk _00866_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[826\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11241__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _02451_ net1538 net238 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05358__Y _01463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11285_ clknet_leaf_63_clk _00797_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[757\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10809__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07854__X _03959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10236_ net1127 net1452 net912 _05226_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_52_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 net1012 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1021 net1024 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1032 net1033 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__buf_4
XFILLER_0_24_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10167_ net123 net916 net906 net1540 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a22o_1
Xfanout1043 net1053 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_4
Xfanout1065 core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_4
X_10098_ net1441 net516 _05158_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__a21o_1
Xfanout1087 net1090 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_4
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09006__B _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06506__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09456__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06646__A _02747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10066__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09022__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06260_ net1059 core.register_file.registers_state\[132\] net688 core.register_file.registers_state\[164\]
+ net660 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__o221a_1
XANTENNA__09208__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05493__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06690__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06191_ net627 _02282_ _02288_ _02295_ net722 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a311o_4
XFILLER_0_114_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08580__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold504 core.register_file.registers_state\[808\] vssd1 vssd1 vccd1 vccd1 net1823
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold515 core.register_file.registers_state\[45\] vssd1 vssd1 vccd1 vccd1 net1834
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 core.register_file.registers_state\[511\] vssd1 vssd1 vccd1 vccd1 net1845
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold537 core.register_file.registers_state\[536\] vssd1 vssd1 vccd1 vccd1 net1856
+ sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap256 _03541_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_1
XFILLER_0_29_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold548 core.register_file.registers_state\[772\] vssd1 vssd1 vccd1 vccd1 net1867
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09950_ net1528 core.CPU_DAT_O\[6\] net798 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
Xhold559 core.register_file.registers_state\[900\] vssd1 vssd1 vccd1 vccd1 net1878
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11734__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08901_ net2331 net370 _04907_ net438 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09881_ net1118 _05067_ net376 net1841 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08195__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload18_A clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__A3 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ net569 net610 net243 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__and3_1
Xhold1204 core.register_file.registers_state\[91\] vssd1 vssd1 vccd1 vccd1 net2523
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06745__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05284__X _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 core.register_file.registers_state\[714\] vssd1 vssd1 vccd1 vccd1 net2534
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06745__B2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05725__A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07416__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1226 core.register_file.registers_state\[473\] vssd1 vssd1 vccd1 vccd1 net2545
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06320__S net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ core.IO_mod.input_reg\[20\] net251 net725 vssd1 vssd1 vccd1 vccd1 _04818_
+ sky130_fd_sc_hd__a21o_1
X_05975_ net1034 core.register_file.registers_state\[717\] core.register_file.registers_state\[749\]
+ net665 net1008 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__o221a_1
XANTENNA__08101__A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05953__C1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ net489 _03721_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09695__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08498__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11269__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ net2011 net467 net434 _04760_ vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__a22o_1
XANTENNA__08595__X _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07645_ _03746_ _03749_ net485 vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07170__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout350_A _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08755__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ _03582_ _03607_ net548 _03680_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08247__S net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06556__A _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09447__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10057__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06527_ _01583_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__xnor2_1
X_09315_ _04939_ net422 net334 net2028 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a22o_1
XANTENNA__09998__B2 _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout236_X net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06458_ net584 _02562_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__or2_1
X_09246_ core.register_file.registers_state\[314\] net474 net544 vssd1 vssd1 vccd1
+ vccd1 _05039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08771__A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06130__C1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05409_ net1059 net754 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_135_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ _04652_ _04660_ _04710_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_135_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06389_ net944 core.register_file.registers_state\[577\] net702 core.register_file.registers_state\[609\]
+ net657 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1145_X net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09214__A3 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ _01365_ _03618_ net547 net504 _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout984_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08059_ net533 _04159_ _04163_ _03685_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__o211a_1
XANTENNA__08973__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1312_X net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ clknet_leaf_93_clk _00582_ net1239 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[542\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net594 _01824_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__nor2_4
XANTENNA__07528__A3 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__A1 core.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05635__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08489__A1 _03536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ clknet_leaf_108_clk _00435_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[395\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07700__A3 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10854_ clknet_leaf_105_clk _00366_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[326\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09438__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07061__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09989__B2 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ clknet_leaf_85_clk _00297_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[257\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07464__A2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09205__A3 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10631__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11406_ clknet_leaf_90_clk _00918_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[878\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07216__A2 _02451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10220__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08964__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11337_ clknet_leaf_16_clk _00849_ net1216 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06975__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11268_ clknet_leaf_75_clk _00780_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[740\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10781__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__A2 _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09913__A1 core.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ net70 net915 vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__and2_1
XANTENNA__06188__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ clknet_leaf_15_clk _00711_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[671\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06727__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05545__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07463__C net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05760_ _01864_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08856__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05691_ net948 core.register_file.registers_state\[821\] net763 net962 vssd1 vssd1
+ vccd1 vccd1 _01796_ sky130_fd_sc_hd__o31a_1
XFILLER_0_72_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07430_ net779 _03528_ _03529_ net767 vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__o31a_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06360__C1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07361_ net969 _03464_ _03465_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06312_ net1062 core.register_file.registers_state\[867\] net754 _02416_ vssd1 vssd1
+ vccd1 vccd1 _02417_ sky130_fd_sc_hd__a31o_1
X_09100_ net2223 net365 net358 _04833_ vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__a22o_1
X_07292_ _03176_ _03205_ _03395_ _03175_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__a31o_2
XANTENNA__07455__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09031_ net742 net462 _04993_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__and3_1
X_06243_ net1059 net755 core.register_file.registers_state\[644\] vssd1 vssd1 vccd1
+ vccd1 _02348_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06174_ net1049 core.register_file.registers_state\[134\] net674 core.register_file.registers_state\[166\]
+ net654 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__o221a_1
XANTENNA__09601__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 core.register_file.registers_state\[545\] vssd1 vssd1 vccd1 vccd1 net1620
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold312 core.register_file.registers_state\[250\] vssd1 vssd1 vccd1 vccd1 net1631
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 net202 vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 core.register_file.registers_state\[261\] vssd1 vssd1 vccd1 vccd1 net1653
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 core.register_file.registers_state\[895\] vssd1 vssd1 vccd1 vccd1 net1664
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 core.register_file.registers_state\[800\] vssd1 vssd1 vccd1 vccd1 net1675
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 core.register_file.registers_state\[825\] vssd1 vssd1 vccd1 vccd1 net1686
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 net102 vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net1010 core.CPU_DAT_O\[22\] net892 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
Xhold389 core.register_file.registers_state\[295\] vssd1 vssd1 vccd1 vccd1 net1708
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_4
XFILLER_0_106_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08168__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout825 net826 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_4
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08707__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout847 net848 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
X_09864_ _04935_ net388 net268 net1839 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout858 net860 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1105_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 core.register_file.registers_state\[589\] vssd1 vssd1 vccd1 vccd1 net2320
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 net871 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05455__A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07146__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1012 core.register_file.registers_state\[100\] vssd1 vssd1 vccd1 vccd1 net2331
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ net462 _04711_ _04862_ net466 net2531 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__a32o_1
Xhold1023 core.register_file.registers_state\[227\] vssd1 vssd1 vccd1 vccd1 net2342
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _04797_ net387 net271 net2197 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__a22o_1
Xhold1034 core.register_file.registers_state\[578\] vssd1 vssd1 vccd1 vccd1 net2353
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06813__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 core.register_file.registers_state\[198\] vssd1 vssd1 vccd1 vccd1 net2364
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1056 core.register_file.registers_state\[862\] vssd1 vssd1 vccd1 vccd1 net2375
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 core.register_file.registers_state\[598\] vssd1 vssd1 vccd1 vccd1 net2386
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ core.IO_mod.data_from_mem\[17\] net246 _04803_ vssd1 vssd1 vccd1 vccd1 _04804_
+ sky130_fd_sc_hd__a21o_2
Xhold1078 core.register_file.registers_state\[843\] vssd1 vssd1 vccd1 vccd1 net2397
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05958_ net1034 core.register_file.registers_state\[461\] core.register_file.registers_state\[493\]
+ net665 net1008 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__o221a_1
XANTENNA__09668__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1089 core.register_file.registers_state\[596\] vssd1 vssd1 vccd1 vccd1 net2408
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08677_ net733 _04172_ _04717_ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__o211a_4
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05889_ net927 _01993_ _01992_ net1029 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__o211a_1
XANTENNA__07143__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1095_X net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07628_ _03655_ _03657_ _03679_ _03690_ _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__a311o_2
XANTENNA__07694__A2 _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07559_ net487 net477 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__nor2_2
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1262_X net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10570_ clknet_leaf_106_clk _00082_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09840__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09229_ _04802_ net417 net339 net1717 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_94_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09199__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10255__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06406__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08946__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09536__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ clknet_leaf_68_clk _00634_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[594\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold890 core.IO_mod.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11053_ clknet_leaf_2_clk _00565_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[525\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10004_ net1465 net540 net519 _05102_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09371__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09659__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06895__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09271__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07580__A _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07134__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906_ clknet_leaf_5_clk _00418_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[378\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07685__A2 _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11886_ clknet_leaf_49_clk _01355_ net1311 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06342__C1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08963__X _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05696__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10837_ clknet_leaf_62_clk _00349_ net1242 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[309\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10755__RESET_B net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09831__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ clknet_leaf_105_clk _00280_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[240\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07739__B _03843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10699_ clknet_leaf_109_clk _00211_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[171\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08937__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06930_ core.register_file.registers_state\[299\] core.register_file.registers_state\[267\]
+ core.register_file.registers_state\[427\] core.register_file.registers_state\[395\]
+ net832 net1069 vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09898__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ _02962_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__and2_1
XANTENNA__06176__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ _03884_ _03964_ _03985_ _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__nand4b_1
X_05812_ net619 _01915_ _01916_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__or3_1
X_06792_ net988 core.register_file.registers_state\[688\] net869 core.register_file.registers_state\[656\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__o221a_1
X_09580_ _04925_ net395 net299 net1789 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08586__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ _04603_ _04604_ _04610_ net208 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a2bb2o_1
X_05743_ core.register_file.registers_state\[20\] net691 net663 _01847_ vssd1 vssd1
+ vccd1 vccd1 _01848_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07125__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_62_clk_X clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10677__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ _04546_ _04547_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__nor2_1
X_05674_ net584 _01747_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07413_ core.register_file.registers_state\[792\] core.register_file.registers_state\[824\]
+ net864 vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__mux2_1
X_08393_ _04483_ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__nor2_1
XANTENNA__06884__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08592__Y _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07344_ _03446_ _03448_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09822__A0 _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05439__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05439__B2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07275_ _03378_ _03379_ net787 vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_132_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06100__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout313_A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1055_A core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09014_ net2437 net427 _04982_ net431 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__a22o_1
X_06226_ _02329_ _02330_ net618 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold1163_A core.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 core.register_file.registers_state\[1\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06157_ core.register_file.registers_state\[935\] core.register_file.registers_state\[903\]
+ net685 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
Xhold131 core.register_file.registers_state\[3\] vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06939__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 net174 vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10196__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__B2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 _01123_ vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11302__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 net178 vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold175 core.IO_mod.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
X_06088_ core.register_file.registers_state\[9\] core.register_file.registers_state\[41\]
+ net699 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold186 core.IO_mod.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout600 _01454_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_2
Xhold197 net197 vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05611__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout611 _04659_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_4
X_09916_ core.control_logic.instruction\[5\] net2483 net891 vssd1 vssd1 vccd1 vccd1
+ _01069_ sky130_fd_sc_hd__mux2_1
Xfanout622 net626 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1010_X net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout633 net635 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_8
Xfanout644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_2
XANTENNA__09889__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1108_X net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 net656 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09353__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _04901_ net390 net268 net1995 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__a22o_1
Xfanout677 net678 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__C_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 net689 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_87_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout947_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05375__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ net562 net458 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_83_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06572__C1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ net728 _04268_ net525 _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_96_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11740_ clknet_leaf_37_clk _01252_ net1223 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06324__C1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11671_ clknet_leaf_36_clk _01183_ net1222 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10622_ clknet_leaf_96_clk _00134_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08616__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09813__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07559__B net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10553_ clknet_leaf_70_clk _00065_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10484_ net1383 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05850__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08919__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09041__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09266__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07052__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__A_N _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05640__A1_N net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ clknet_leaf_101_clk _00617_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[577\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09344__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ clknet_leaf_42_clk _00548_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[508\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06563__C1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07107__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08693__X _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05669__A1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11869_ clknet_leaf_52_clk _01338_ net1303 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06961__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05390_ net1123 _01404_ _01492_ _01494_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__and4_2
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09804__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09030__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06618__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09280__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07060_ net974 _03161_ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a21o_1
XANTENNA__11325__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06011_ core.decoder.inst\[7\] _01387_ _01402_ _01391_ net1052 vssd1 vssd1 vccd1
+ vccd1 _02116_ sky130_fd_sc_hd__a32o_1
XANTENNA__05841__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05841__B2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10178__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07043__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08240__C1 _02488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09583__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06397__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07962_ _02084_ _02931_ _03621_ _02053_ net900 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__a32o_1
XANTENNA__07772__X _03877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _04891_ net2044 net281 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06913_ net1098 core.register_file.registers_state\[332\] core.register_file.registers_state\[364\]
+ net841 net980 vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07893_ net1003 _03996_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08587__Y _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09632_ net745 _05005_ net459 vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and3_1
X_06844_ net777 _02945_ _02948_ net773 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__a31o_1
XANTENNA__10350__A0 _05102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07897__A2 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09563_ net203 net2431 net303 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__mux2_1
X_06775_ net784 _02878_ _02879_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _01384_ _03475_ net574 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__mux2_1
X_05726_ net1065 core.register_file.registers_state\[852\] vssd1 vssd1 vccd1 vccd1
+ _01831_ sky130_fd_sc_hd__or2_1
X_09494_ net603 net203 net319 net261 net1745 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__a32o_1
X_08445_ _01828_ _04530_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05657_ _01753_ _01756_ _01758_ _01761_ net934 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_114_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_42_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1172_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08059__C1 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08376_ core.pc.current_pc\[14\] _02994_ net576 vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__mux2_1
X_05588_ net1011 _01690_ _01691_ net959 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_119_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07327_ net969 _03423_ _03431_ net775 vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a211o_1
XANTENNA__09271__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09810__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07258_ net996 core.register_file.registers_state\[960\] net888 core.register_file.registers_state\[992\]
+ net977 vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06209_ _02296_ _02313_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__nand2_8
X_07189_ core.register_file.registers_state\[802\] core.register_file.registers_state\[770\]
+ core.register_file.registers_state\[930\] core.register_file.registers_state\[898\]
+ net854 net1078 vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09023__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10169__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09574__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07585__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08782__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__X _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06793__C1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _04962_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_8
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_2
XANTENNA__10842__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout452 net454 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_2
XANTENNA__09326__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09814__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 net465 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07337__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout485 _02516_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07337__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout496 _02486_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09877__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05348__B1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10341__A0 _02421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05899__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10992__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11723_ clknet_leaf_48_clk _01235_ net1306 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ clknet_leaf_47_clk _01166_ net1306 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08018__X _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06474__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10605_ clknet_leaf_0_clk _00117_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09262__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ clknet_leaf_27_clk _01097_ net1197 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09801__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07273__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10536_ clknet_leaf_95_clk _00048_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05823__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05284__C1 core.decoder.inst\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ net1382 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09014__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07576__A1 _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ net1391 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07120__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09009__B _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__X _03697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09317__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08848__B _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ clknet_leaf_111_clk _00531_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[491\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10332__A0 _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__Y _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09025__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05272__B core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ core.register_file.registers_state\[791\] core.register_file.registers_state\[823\]
+ core.register_file.registers_state\[919\] core.register_file.registers_state\[951\]
+ net866 net1071 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05511_ _01500_ _01615_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__nor2_1
XANTENNA__06839__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06491_ net631 _02592_ _02595_ net721 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09679__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07500__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ _01495_ _03740_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__nor2_4
X_05442_ net963 _01543_ net629 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09398__C net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10715__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08161_ net265 _04159_ _04168_ _04024_ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__a221o_1
X_05373_ net1100 core.register_file.registers_state\[990\] core.register_file.registers_state\[1022\]
+ net843 net1075 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06067__A1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ _03212_ _03215_ _03216_ _03209_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__o22a_1
X_08092_ net495 _04147_ _04196_ net534 vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload40 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_12
X_07043_ net1107 core.register_file.registers_state\[135\] net848 core.register_file.registers_state\[167\]
+ net824 vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload51 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_110_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__B _01987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload62 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_8
Xclkload73 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_8
XANTENNA__09005__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__inv_6
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload95 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ net614 net223 vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1018_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09308__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ _02146_ _03052_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__and2_1
XANTENNA__07319__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07319__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07876_ net531 _03696_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05463__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07154__S net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09615_ net2151 net391 _05070_ net998 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06827_ net538 _02526_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout645_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09546_ net206 net2289 net306 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__mux2_1
X_06758_ core.register_file.registers_state\[721\] core.register_file.registers_state\[753\]
+ net883 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__mux2_1
XANTENNA__08774__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05709_ net1056 core.register_file.registers_state\[181\] vssd1 vssd1 vccd1 vccd1
+ _01814_ sky130_fd_sc_hd__and2_1
X_09477_ _04985_ net318 net262 net1905 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout812_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06689_ core.register_file.registers_state\[531\] core.register_file.registers_state\[563\]
+ net869 vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09492__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05728__S1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08428_ _04515_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_117_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06294__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05502__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload1 clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ _04431_ _04435_ _04445_ _04443_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o31a_1
XFILLER_0_74_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11370_ clknet_leaf_111_clk _00882_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[842\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05805__A1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05805__B2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10321_ _05106_ net1483 net237 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
X_10252_ net1125 net1478 net910 _05234_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__a31o_1
XANTENNA__11790__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06233__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ net110 net918 net908 net1485 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a22o_1
XANTENNA__05357__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1203 net1208 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05569__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1214 net1216 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_4
Xfanout1225 net1226 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09544__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06230__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05664__S0 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1236 net1250 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_2
XANTENNA_input39_A gpio_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1247 net1249 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__clkbuf_4
Xfanout260 _05084_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_4
Xfanout1258 net1262 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1269 net1271 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_4
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
XANTENNA__10314__A0 _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout293 net298 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09180__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07191__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11170__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08684__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05741__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10738__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09499__B net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09483__A1 _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06297__A1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ clknet_leaf_52_clk net1534 net1302 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08691__C1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11637_ clknet_leaf_53_clk _01149_ net1302 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09235__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06049__A1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09786__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08589__A3 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ clknet_leaf_28_clk _01080_ net1194 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07797__A1 core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold708 core.register_file.registers_state\[665\] vssd1 vssd1 vccd1 vccd1 net2027
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ clknet_leaf_35_clk _00031_ net1219 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold719 core.register_file.registers_state\[41\] vssd1 vssd1 vccd1 vccd1 net2038
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11499_ clknet_leaf_110_clk _01011_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[971\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06221__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05991_ net655 _02090_ _02091_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__o21a_1
XANTENNA__08578__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ net495 _03654_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__nor2_1
XANTENNA__10305__A0 _02451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05980__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06509__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10897__Q core.register_file.registers_state\[369\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09171__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07661_ net500 net454 _03231_ net446 vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07721__B2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ net2253 net226 net407 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06612_ net769 _02711_ _02716_ _02704_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a31o_4
X_07592_ _02385_ _03656_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__or2_4
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08594__A core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10069__C1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09331_ net464 _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__nand2_1
X_06543_ net1104 core.register_file.registers_state\[988\] core.register_file.registers_state\[1020\]
+ net852 net1077 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08277__A2 _01412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06288__A1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ net2302 net225 net338 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06474_ net1004 _02577_ _02578_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08213_ _03964_ _04278_ _04286_ _04306_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__and4b_1
XANTENNA__05496__C1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05425_ net962 _01529_ _01528_ net1017 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a211o_1
X_09193_ _04991_ net357 net425 net1765 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout226_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08144_ net1113 _02385_ _03261_ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__o31a_1
X_05356_ core.register_file.registers_state\[30\] core.register_file.registers_state\[62\]
+ core.register_file.registers_state\[158\] core.register_file.registers_state\[190\]
+ net870 net820 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__mux4_1
XANTENNA__09777__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08075_ _03797_ _03858_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05287_ _01364_ _01401_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__and2_1
XANTENNA__06996__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1135_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06460__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07026_ net1101 core.register_file.registers_state\[584\] core.register_file.registers_state\[616\]
+ net845 net807 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__o221a_1
XANTENNA__05458__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1302_A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06212__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 core.register_file.registers_state\[19\] vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 core.register_file.registers_state\[9\] vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ net243 net736 vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__and2_1
Xhold35 core.register_file.registers_state\[980\] vssd1 vssd1 vccd1 vccd1 net1354
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_A _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 core.register_file.registers_state\[952\] vssd1 vssd1 vccd1 vccd1 net1365
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _01987_ _02873_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__or2_1
Xhold57 core.register_file.registers_state\[1020\] vssd1 vssd1 vccd1 vccd1 net1376
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 core.register_file.registers_state\[978\] vssd1 vssd1 vccd1 vccd1 net1387
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11193__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold79 core.register_file.registers_state\[999\] vssd1 vssd1 vccd1 vccd1 net1398
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _03548_ net529 _03947_ _03963_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout1292_X net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05723__B1 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ clknet_leaf_43_clk _00382_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ _04867_ net403 net310 net1869 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06279__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09217__A1 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08951__B _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09539__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11422_ clknet_leaf_95_clk _00934_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[894\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07779__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ clknet_leaf_64_clk _00865_ net1267 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06987__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10304_ _04229_ net245 vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__nand2b_1
XANTENNA__05368__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06451__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05885__S0 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11284_ clknet_leaf_51_clk _00796_ net1297 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[756\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10235_ net78 net915 vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06898__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08679__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1000 net1002 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_4
XANTENNA__11536__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09274__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_37_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1022 net1024 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_37_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1033 core.decoder.inst\[21\] vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_6
X_10166_ net112 net916 net906 net1512 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a22o_1
Xfanout1044 net1050 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
Xfanout1055 core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_8
Xfanout1077 net1081 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_4
X_10097_ _04298_ net557 net588 core.pc.current_pc\[18\] net471 vssd1 vssd1 vccd1 vccd1
+ _05158_ sky130_fd_sc_hd__o221a_1
XANTENNA__06199__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_4
XFILLER_0_89_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1099 net1103 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
XANTENNA__09153__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07703__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06911__C1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10999_ clknet_leaf_22_clk _00511_ net1181 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[471\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06190_ net960 _02289_ _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09759__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06690__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold505 core.register_file.registers_state\[277\] vssd1 vssd1 vccd1 vccd1 net1824
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 core.register_file.registers_state\[817\] vssd1 vssd1 vccd1 vccd1 net1835
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 core.register_file.registers_state\[492\] vssd1 vssd1 vccd1 vccd1 net1846
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 core.register_file.registers_state\[565\] vssd1 vssd1 vccd1 vccd1 net1857
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 core.register_file.registers_state\[57\] vssd1 vssd1 vccd1 vccd1 net1868
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ net572 net223 net737 vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__and3_2
XFILLER_0_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09880_ net1119 _04964_ net461 net377 net1554 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08195__A1 _01781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08195__B2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07493__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ net607 _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1205 core.register_file.registers_state\[337\] vssd1 vssd1 vccd1 vccd1 net2524
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05548__A3 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1216 core.register_file.registers_state\[183\] vssd1 vssd1 vccd1 vccd1 net2535
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10903__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ net1904 net466 net433 _04817_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__a22o_1
Xhold1227 core.register_file.registers_state\[369\] vssd1 vssd1 vccd1 vccd1 net2546
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05974_ net1034 core.register_file.registers_state\[589\] core.register_file.registers_state\[621\]
+ net665 net923 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07713_ net512 _03817_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__nor2_1
XANTENNA__09912__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ net567 _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__and2_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07644_ _03747_ _03748_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08755__C net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07575_ net1114 _03608_ net580 core.decoder.inst\[31\] net899 vssd1 vssd1 vccd1 vccd1
+ _03680_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout343_A _05027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ net559 _04937_ _05049_ net331 net2440 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06526_ _01612_ _02601_ net537 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__o21a_1
XANTENNA__09998__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__B net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11238__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05469__C1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09500__X _05063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09245_ net561 _04851_ _05038_ net342 net2538 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout510_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06457_ core.decoder.inst\[24\] net899 net593 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__B _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1252_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07668__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05408_ net940 net761 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__nor2_1
X_09176_ net242 net739 net358 net345 net2047 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_135_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06388_ core.register_file.registers_state\[545\] core.register_file.registers_state\[513\]
+ net682 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08127_ net497 _04231_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05339_ net1129 net1911 _01423_ _01427_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08058_ net533 _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_92_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_A _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ _02206_ _03113_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__xor2_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1305_X net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07607__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ net1572 net541 net520 _05110_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__a22o_1
XANTENNA__06197__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__A1 _04037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__D1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__X _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05944__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09822__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10922_ clknet_leaf_106_clk _00434_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[394\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06747__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11899__1316 vssd1 vssd1 vccd1 vccd1 _11899__1316/HI net1316 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_45_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10853_ clknet_leaf_87_clk _00365_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[325\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05370__B net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ clknet_leaf_55_clk _00296_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[256\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08962__A _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09269__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06672__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ clknet_leaf_0_clk _00917_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[877\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05880__C1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07621__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11336_ clknet_leaf_9_clk _00848_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08612__D_N _03964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07584__Y _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ clknet_leaf_67_clk _00779_ net1268 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[739\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08177__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__B1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ net1127 net1509 net912 _05217_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__a31o_1
X_11198_ clknet_leaf_95_clk _00710_ net1178 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[670\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07385__C1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10149_ net470 _05195_ _05197_ net515 net1484 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a32o_1
XANTENNA__09126__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05935__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07137__C1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__B _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05690_ net948 core.register_file.registers_state\[885\] net763 _01791_ net1029 vssd1
+ vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__o311a_1
XANTENNA__07252__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09033__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05699__C1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire409_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09429__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06360__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05280__B core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07360_ net1094 core.register_file.registers_state\[858\] core.register_file.registers_state\[890\]
+ net836 net978 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08872__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06311_ net954 core.register_file.registers_state\[835\] net1020 vssd1 vssd1 vccd1
+ vccd1 _02416_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07291_ _03205_ _03395_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__and2_1
XANTENNA__06112__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09030_ net612 net218 vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06242_ core.decoder.inst\[11\] _01409_ _01411_ core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 _02347_ sky130_fd_sc_hd__a22oi_4
XANTENNA__06663__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05466__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06663__B2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05871__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06173_ net585 _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__nor2_1
Xhold302 net159 vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09601__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 core.i_hit vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06415__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold324 core.register_file.registers_state\[389\] vssd1 vssd1 vccd1 vccd1 net1643
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold335 core.register_file.registers_state\[810\] vssd1 vssd1 vccd1 vccd1 net1654
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold346 core.register_file.registers_state\[390\] vssd1 vssd1 vccd1 vccd1 net1665
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 core.register_file.registers_state\[543\] vssd1 vssd1 vccd1 vccd1 net1676
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net1026 core.CPU_DAT_O\[21\] net894 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold368 core.register_file.registers_state\[386\] vssd1 vssd1 vccd1 vccd1 net1687
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold379 net200 vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout804 net807 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout815 _01460_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout826 _01459_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_4
XANTENNA__05736__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout837 net838 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_4
X_09863_ net561 _04933_ net459 net267 net1684 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout293_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_2
Xhold1002 core.register_file.registers_state\[328\] vssd1 vssd1 vccd1 vccd1 net2321
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08814_ net565 _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and2_1
Xhold1013 core.register_file.registers_state\[88\] vssd1 vssd1 vccd1 vccd1 net2332
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09794_ net569 _04791_ net387 net271 net1674 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__a32o_1
Xhold1024 core.register_file.registers_state\[622\] vssd1 vssd1 vccd1 vccd1 net2343
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 core.register_file.registers_state\[65\] vssd1 vssd1 vccd1 vccd1 net2354
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06194__A3 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1046 core.register_file.registers_state\[851\] vssd1 vssd1 vccd1 vccd1 net2365
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ core.IO_mod.input_reg\[17\] net250 net725 vssd1 vssd1 vccd1 vccd1 _04803_
+ sky130_fd_sc_hd__a21o_1
Xhold1057 core.register_file.registers_state\[220\] vssd1 vssd1 vccd1 vccd1 net2376
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 core.register_file.registers_state\[832\] vssd1 vssd1 vccd1 vccd1 net2387
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05957_ net1036 core.register_file.registers_state\[333\] core.register_file.registers_state\[365\]
+ net665 net923 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout460_A _05060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 core.register_file.registers_state\[880\] vssd1 vssd1 vccd1 vccd1 net2398
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08766__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10278__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ core.IO_mod.data_from_mem\[6\] net247 _04744_ vssd1 vssd1 vccd1 vccd1 _04745_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05888_ net946 core.register_file.registers_state\[463\] net704 core.register_file.registers_state\[495\]
+ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
XANTENNA__06567__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _03697_ _03731_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout725_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1088_X net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ net498 net451 _02660_ net443 vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06509_ net1096 core.register_file.registers_state\[477\] core.register_file.registers_state\[509\]
+ net837 net1070 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07489_ net967 _03589_ _03592_ _03593_ _03584_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09228_ _04797_ net421 net341 net2035 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__a22o_1
XANTENNA__05457__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09159_ _04926_ net357 net345 net2080 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06406__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09817__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ clknet_leaf_74_clk _00633_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[593\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08159__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold880 core.register_file.registers_state\[477\] vssd1 vssd1 vccd1 vccd1 net2199
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold891 core.register_file.registers_state\[170\] vssd1 vssd1 vccd1 vccd1 net2210
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09356__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05646__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ clknet_leaf_102_clk _00564_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[524\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07367__C1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ net724 _02113_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__and2_2
XFILLER_0_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05917__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__RESET_B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06017__S0 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07072__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10905_ clknet_leaf_55_clk _00417_ net1295 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[377\]
+ sky130_fd_sc_hd__dfrtp_1
X_11885_ clknet_leaf_47_clk _01354_ net1292 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06342__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05696__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10836_ clknet_leaf_56_clk _00348_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[308\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08692__A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10767_ clknet_leaf_82_clk _00279_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[239\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06924__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ clknet_leaf_106_clk _00210_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09595__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06948__A2 _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07896__A2_N _03843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11319_ clknet_leaf_7_clk _00831_ net1182 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[791\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap523_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09347__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09028__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09898__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06860_ _02016_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__xnor2_1
X_05811_ net1060 core.register_file.registers_state\[210\] core.register_file.registers_state\[242\]
+ net690 net662 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__o221a_1
X_06791_ core.register_file.registers_state\[528\] core.register_file.registers_state\[560\]
+ net869 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__mux2_1
XANTENNA__08586__B net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ _04605_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05742_ net1063 core.register_file.registers_state\[52\] net755 vssd1 vssd1 vccd1
+ vccd1 _01847_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08322__A1 _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08461_ _01782_ _04543_ _04544_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05673_ _01764_ _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07412_ _03513_ _03514_ _03516_ _03515_ net789 net802 vssd1 vssd1 vccd1 vccd1 _03517_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06884__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ _01988_ _04481_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07343_ _01708_ _03447_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06097__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09985__X _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09210__B _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06636__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07274_ net996 core.register_file.registers_state\[192\] net889 core.register_file.registers_state\[224\]
+ net814 vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_14_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06636__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09013_ net563 _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__and2_1
XANTENNA__05844__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06225_ net944 core.register_file.registers_state\[709\] net702 core.register_file.registers_state\[741\]
+ net643 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08389__A1 _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1048_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold110 core.register_file.registers_state\[984\] vssd1 vssd1 vccd1 vccd1 net1429
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09586__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 core.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ net948 core.register_file.registers_state\[839\] net706 core.register_file.registers_state\[871\]
+ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a22o_1
Xhold132 core.IO_mod.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09050__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 core.register_file.registers_state\[18\] vssd1 vssd1 vccd1 vccd1 net1462
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 core.ru.state\[1\] vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold165 core.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06087_ core.register_file.registers_state\[201\] core.register_file.registers_state\[233\]
+ net699 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
Xhold176 core.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1215_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 net158 vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _04897_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_4
XANTENNA__09338__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold198 core.CPU_DAT_I\[4\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05611__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout612 net615 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_4
X_09915_ net1123 core.CPU_DAT_O\[4\] net893 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__mux2_1
Xfanout623 net625 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
XFILLER_0_10_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07349__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout675_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 net650 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout656 net664 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_4
X_09846_ _04899_ net388 net267 net2330 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__a22o_1
Xfanout667 net680 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__A core.IO_mod.input_reg\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_87_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 _01514_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_87_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05375__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ _05020_ net290 net259 net2235 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__a22o_1
X_06989_ net1085 _03093_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08728_ core.IO_mod.data_from_mem\[14\] net249 _04788_ vssd1 vssd1 vccd1 vccd1 _04789_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__05913__B _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10311__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10621__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11253__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09510__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08659_ net609 net224 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06324__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ clknet_leaf_36_clk _01182_ net1222 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ clknet_leaf_17_clk _00133_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08616__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07824__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10552_ clknet_leaf_10_clk _00064_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10483_ net1345 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11127__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09577__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09547__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09041__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07052__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06486__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11104_ clknet_leaf_58_clk _00616_ net1287 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[576\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06260__C1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09329__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11277__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05807__C net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ clknet_leaf_19_clk _00547_ net1191 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[507\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07591__A _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05366__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05366__B2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06563__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09501__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08599__A_N _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05542__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11868_ clknet_leaf_53_clk _01337_ net1300 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06961__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10819_ clknet_leaf_73_clk _00331_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11799_ clknet_leaf_50_clk _01300_ net1307 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09804__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06079__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09030__B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05826__C1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06010_ _01408_ _01424_ core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__o21a_1
XANTENNA__05985__S net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09568__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09032__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07043__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07594__A2 _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ _02937_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09700_ net214 net2184 net281 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
X_06912_ core.register_file.registers_state\[268\] core.register_file.registers_state\[300\]
+ core.register_file.registers_state\[396\] core.register_file.registers_state\[428\]
+ net870 net1073 vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07892_ net1032 net900 net548 _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a22o_1
XANTENNA__08543__A1 _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ _05004_ net399 net393 net1881 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__a22o_1
X_06843_ _02946_ _02947_ net786 vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ net210 net2486 net305 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06774_ net1093 core.register_file.registers_state\[208\] core.register_file.registers_state\[240\]
+ net833 net817 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__o221a_1
XANTENNA__09099__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ net208 _04592_ _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__or3_1
XANTENNA__09920__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05725_ net955 core.register_file.registers_state\[884\] net766 vssd1 vssd1 vccd1
+ vccd1 _01830_ sky130_fd_sc_hd__or3_1
XANTENNA__10794__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06306__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ _05015_ net322 net264 net1626 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a22o_1
X_08444_ _01828_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06857__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05656_ net659 _01759_ _01760_ net1030 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08375_ net2551 _04468_ net599 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__mux2_1
X_05587_ net1042 core.register_file.registers_state\[347\] core.register_file.registers_state\[379\]
+ net671 net922 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout423_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06609__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07326_ _03424_ _03425_ net1090 vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__o21a_1
XANTENNA__10646__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06609__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06056__S net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10086__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07257_ core.register_file.registers_state\[800\] core.register_file.registers_state\[768\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11499__SET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06208_ net717 _02303_ _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__or3b_4
XFILLER_0_131_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08124__X _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07188_ _03289_ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nand2_1
XANTENNA__09023__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07034__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06139_ core.register_file.registers_state\[167\] net681 net657 _02243_ vssd1 vssd1
+ vccd1 vccd1 _02244_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10306__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1120_X net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07585__A2 _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 net422 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
XANTENNA__05627__C net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 net432 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_4
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 _03630_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_8
Xfanout475 _04666_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout486 _02516_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09731__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout497 net499 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_2
X_09829_ _04800_ net2430 net382 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06298__Y _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09830__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08954__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11722_ clknet_leaf_36_clk _01234_ net1219 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06312__A3 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07350__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ clknet_leaf_36_clk _01165_ net1219 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ clknet_leaf_101_clk _00116_ net1162 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09798__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ clknet_3_2_0_clk _01096_ net1204 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10517__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07273__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10535_ clknet_leaf_91_clk _00047_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05284__B1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09277__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05823__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10466_ net1410 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09014__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07025__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07025__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ net1578 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10667__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07120__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05587__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05587__B2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05393__X _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09722__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ clknet_leaf_0_clk _00530_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11104__RESET_B net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09025__B net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05272__C core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05510_ _01400_ _01614_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__or2_1
XANTENNA__06839__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06490_ _02593_ _02594_ net1025 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08209__X _04314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06303__A3 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05441_ _01544_ _01545_ net1027 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ _03791_ _04018_ _04262_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_clk_X clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09789__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05372_ net1086 _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__or2_1
XANTENNA__09253__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07111_ net1086 _03206_ _03207_ net967 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08091_ net486 _04182_ _04195_ net490 vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload30 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_6
X_07042_ _03052_ _03055_ _03145_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__a211o_1
Xclkload41 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06472__C1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload52 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__inv_6
XANTENNA__09005__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__C _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload63 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__inv_8
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_clk_X clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload74 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_110_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload85 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__inv_6
XANTENNA__09982__Y _05093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload96 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_6
XANTENNA__11592__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10020__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06224__C1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ net2265 net430 _04968_ net1001 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__a22o_1
X_07944_ _03971_ _04015_ net495 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__mux2_2
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ net510 _03697_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_108_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_A _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09614_ net742 _04983_ net456 vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__and3_1
X_06826_ net771 _02917_ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a21o_4
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09545_ net222 net2149 net303 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10898__RESET_B net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06757_ core.register_file.registers_state\[657\] core.register_file.registers_state\[689\]
+ net883 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout638_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05708_ core.register_file.registers_state\[21\] net684 net659 _01812_ vssd1 vssd1
+ vccd1 vccd1 _01813_ sky130_fd_sc_hd__a211o_1
X_09476_ _04983_ net315 net261 net1747 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06688_ net971 _02791_ _02792_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__or3_1
XANTENNA__09492__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08427_ _04512_ _04514_ net229 vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_114_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05639_ net632 _01740_ _01743_ net722 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a31o_1
XANTENNA__05502__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08358_ _04451_ _04452_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__nor2_1
Xclkload2 clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__inv_12
XANTENNA__09244__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07309_ _02717_ _02719_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__and2_1
XANTENNA__07255__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06058__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08452__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ _04366_ _04368_ _04378_ _04380_ _04388_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__o311a_1
XFILLER_0_22_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06581__Y _02686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10320_ _05105_ net1514 net236 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ net87 net914 vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__and2_1
XANTENNA__09952__A0 core.IO_mod.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ net109 net918 net908 net1533 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1208 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1215 net1216 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__clkbuf_4
Xfanout1226 net1236 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05664__S1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1237 net1239 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_4
Xfanout250 net252 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08301__Y _04401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_4
Xfanout1259 net1262 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_50_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_8
Xfanout283 _05081_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_4
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_4
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07191__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__A _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09560__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05741__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08684__B _04751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09483__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07080__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11465__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ clknet_leaf_70_clk net1591 net1275 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07494__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11636_ clknet_leaf_70_clk _01148_ net1274 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09235__A2 _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11567_ clknet_leaf_24_clk _01079_ net1185 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08589__A4 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07797__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10518_ clknet_leaf_36_clk _00030_ net1219 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold709 core.register_file.registers_state\[372\] vssd1 vssd1 vccd1 vccd1 net2028
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ clknet_leaf_111_clk _01010_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[970\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11482__SET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10449_ net1381 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06206__C1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_41_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05990_ net654 _02093_ _02094_ _02092_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09036__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06012__X _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05980__A1 core.decoder.inst\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__inv_2
XANTENNA__06947__X _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05851__X _01956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ net976 _02712_ _02715_ net777 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10991__RESET_B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07591_ _02385_ _03656_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__nor2_1
XANTENNA__08594__B _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10069__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09330_ net1118 net743 net614 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__and3_1
X_06542_ core.register_file.registers_state\[796\] core.register_file.registers_state\[828\]
+ core.register_file.registers_state\[924\] core.register_file.registers_state\[956\]
+ net881 net1077 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09474__A2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ net2131 net227 net337 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06473_ net1034 core.register_file.registers_state\[600\] core.register_file.registers_state\[632\]
+ net666 net636 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08212_ net529 _04307_ _04308_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a31o_2
XANTENNA__07778__X _03883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05424_ core.register_file.registers_state\[798\] core.register_file.registers_state\[830\]
+ net707 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__mux2_1
X_09192_ _04989_ net357 net425 net1727 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload60_A clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ _02385_ _03261_ _03618_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07237__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05355_ _01387_ _01389_ _01392_ _01394_ net979 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a221o_4
XFILLER_0_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload107_A clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06445__C1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _03618_ _04177_ _04178_ net546 _04176_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__o32a_1
XFILLER_0_114_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05286_ core.control_logic.instruction\[2\] core.control_logic.instruction\[0\] core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__and3b_1
XANTENNA__05799__A1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07025_ net1101 core.register_file.registers_state\[712\] core.register_file.registers_state\[744\]
+ net845 net821 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__o221a_1
XANTENNA__06460__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1128_A _01379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__A0 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A _05093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold14 core.register_file.registers_state\[949\] vssd1 vssd1 vccd1 vccd1 net1333
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ net2466 net367 _04957_ net432 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__a22o_1
XANTENNA__11338__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold25 core.register_file.registers_state\[937\] vssd1 vssd1 vccd1 vccd1 net1344
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05420__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 core.register_file.registers_state\[981\] vssd1 vssd1 vccd1 vccd1 net1355
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 core.register_file.registers_state\[8\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ net1003 _01987_ _02873_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nand3_1
Xhold58 core.register_file.registers_state\[964\] vssd1 vssd1 vccd1 vccd1 net1377
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 core.register_file.registers_state\[976\] vssd1 vssd1 vccd1 vccd1 net1388
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05971__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05971__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout755_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__S1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _03696_ _03951_ _03958_ _03962_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__a211o_2
XANTENNA__06857__X _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ net1092 core.register_file.registers_state\[973\] core.register_file.registers_state\[1005\]
+ net831 vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05723__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ net497 _03671_ _03806_ net482 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout922_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05480__Y _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ _04711_ _04862_ net456 net307 net2501 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06279__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ _04952_ net317 net311 net1933 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06684__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09217__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11421_ clknet_leaf_18_clk _00933_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[893\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07228__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08976__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05649__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11352_ clknet_leaf_3_clk _00864_ net1150 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[824\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10303_ _01426_ _04242_ _04695_ _04697_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__nor4_1
XFILLER_0_120_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05885__S1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11283_ clknet_leaf_11_clk _00795_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[755\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08728__A1 core.IO_mod.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__A0 core.decoder.inst\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ net1126 net1441 net912 _05225_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__a31o_1
XANTENNA_input51_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08679__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
Xfanout1012 net1016 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__buf_2
X_10165_ net101 net918 net908 net1804 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__a22o_1
XANTENNA__07583__B _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05384__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07075__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1045 net1050 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_2
Xfanout1056 net1057 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_2
X_10096_ net1425 net518 _05157_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__a21o_1
Xfanout1067 core.decoder.inst\[18\] vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
Xfanout1089 net1090 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07164__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09290__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10855__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ clknet_leaf_44_clk _00510_ net1286 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[470\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09456__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07104__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07011__S0 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07467__B2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09208__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11619_ clknet_leaf_31_clk _01131_ net1201 vssd1 vssd1 vccd1 vccd1 core.WRITE_I sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08967__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold506 core.register_file.registers_state\[888\] vssd1 vssd1 vccd1 vccd1 net1825
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold517 core.register_file.registers_state\[919\] vssd1 vssd1 vccd1 vccd1 net1836
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 core.register_file.registers_state\[63\] vssd1 vssd1 vccd1 vccd1 net1847
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 core.register_file.registers_state\[794\] vssd1 vssd1 vccd1 vccd1 net1858
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09916__A0 core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09465__S net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08195__A2 _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ net727 _04873_ _04874_ net526 vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__o211a_4
Xhold1206 core.register_file.registers_state\[739\] vssd1 vssd1 vccd1 vccd1 net2525
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ net563 net606 net215 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__and3_2
Xhold1217 core.register_file.registers_state\[343\] vssd1 vssd1 vccd1 vccd1 net2536
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05725__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1228 core.register_file.registers_state\[74\] vssd1 vssd1 vccd1 vccd1 net2547
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05973_ net1008 _02077_ _02076_ net932 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a211o_1
XANTENNA__05953__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05953__B2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ _03705_ _03729_ net489 vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__mux2_2
X_08692_ _04670_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07643_ net452 _03052_ net444 net509 vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07574_ net489 _03678_ _03669_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11780__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09447__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09313_ core.register_file.registers_state\[371\] net474 net544 vssd1 vssd1 vccd1
+ vccd1 _05049_ sky130_fd_sc_hd__o21a_1
X_06525_ net767 _02629_ _02617_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__o21a_4
XANTENNA__07014__A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout336_A _05046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09244_ core.register_file.registers_state\[313\] net475 net545 vssd1 vssd1 vccd1
+ vccd1 _05038_ sky130_fd_sc_hd__o21a_1
XANTENNA__06666__C1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06456_ _02535_ _02560_ net584 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__mux2_4
XFILLER_0_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06130__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05407_ core.decoder.inst\[24\] net748 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__nand2_1
XANTENNA__11010__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09175_ _04958_ net354 net344 net2115 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07668__B _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06387_ core.register_file.registers_state\[801\] core.register_file.registers_state\[769\]
+ core.register_file.registers_state\[929\] core.register_file.registers_state\[897\]
+ net682 net1017 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_135_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11278__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ net579 net530 vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nor2_1
X_05338_ net1315 _01427_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_96_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08958__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07955__Y _04060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08057_ _04081_ _04099_ _04138_ _04160_ net478 net494 vssd1 vssd1 vccd1 vccd1 _04162_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07091__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05269_ core.pc.current_pc\[26\] vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06999__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07008_ _02241_ _02524_ net539 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09907__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10728__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06197__A1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ net212 net735 vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_32_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10921_ clknet_leaf_16_clk _00433_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[393\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10852_ clknet_leaf_75_clk _00364_ net1262 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[324\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09438__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10783_ clknet_leaf_94_clk _00295_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[255\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08962__B net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08110__A2 _04100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06121__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08949__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ clknet_leaf_103_clk _00916_ net1156 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09071__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09610__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11335_ clknet_leaf_65_clk _00847_ net1246 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[807\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10220__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ clknet_leaf_78_clk _00778_ net1253 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[738\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10217_ net69 net915 vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__and2_1
XANTENNA__11653__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06188__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ clknet_leaf_20_clk _00709_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[669\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10148_ net556 _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nand2_1
XANTENNA__06003__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05545__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08696__Y _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10079_ _04064_ net590 vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__nand2_1
XANTENNA__09677__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09033__B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06360__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11033__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08872__B _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06310_ net1054 core.register_file.registers_state\[995\] net753 _02414_ net929 vssd1
+ vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a311o_1
XFILLER_0_58_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07769__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__C1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07290_ _03236_ _03393_ _03204_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a21o_1
XANTENNA__06112__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06241_ net582 _02343_ _02344_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_127_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11371__RESET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05289__A core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06172_ core.decoder.inst\[26\] net734 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold303 core.register_file.registers_state\[791\] vssd1 vssd1 vccd1 vccd1 net1622
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 core.register_file.registers_state\[779\] vssd1 vssd1 vccd1 vccd1 net1633
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06415__A2 _02381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 core.register_file.registers_state\[287\] vssd1 vssd1 vccd1 vccd1 net1644
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold336 core.ADR_I\[5\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 core.IO_mod.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold358 core.register_file.registers_state\[293\] vssd1 vssd1 vccd1 vccd1 net1677
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05623__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09931_ net1042 net2553 net894 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
Xhold369 core.register_file.registers_state\[746\] vssd1 vssd1 vccd1 vccd1 net1688
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06820__C1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
Xfanout816 net818 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_4
X_09862_ _04931_ net385 net269 net2398 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__a22o_1
XANTENNA__06179__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout827 net830 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_4
XANTENNA__09904__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout838 _01458_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08887__X _04898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout849 net861 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07915__A2 _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07009__A _02206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ net605 _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__nor2_1
Xhold1003 core.register_file.registers_state\[70\] vssd1 vssd1 vccd1 vccd1 net2322
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 core.register_file.registers_state\[347\] vssd1 vssd1 vccd1 vccd1 net2333
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _04787_ net383 net270 net1988 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1025 core.register_file.registers_state\[920\] vssd1 vssd1 vccd1 vccd1 net2344
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 core.register_file.registers_state\[732\] vssd1 vssd1 vccd1 vccd1 net2355
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 core.register_file.registers_state\[62\] vssd1 vssd1 vccd1 vccd1 net2366
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ net1970 net466 net432 _04802_ vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__a22o_1
X_05956_ core.register_file.registers_state\[269\] core.register_file.registers_state\[301\]
+ core.register_file.registers_state\[397\] core.register_file.registers_state\[429\]
+ net695 net1009 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__mux4_1
Xhold1058 core.register_file.registers_state\[840\] vssd1 vssd1 vccd1 vccd1 net2377
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 core.register_file.registers_state\[157\] vssd1 vssd1 vccd1 vccd1 net2388
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09668__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ core.IO_mod.input_reg\[6\] net251 net726 vssd1 vssd1 vccd1 vccd1 _04744_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__07679__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05887_ net946 core.register_file.registers_state\[335\] net704 core.register_file.registers_state\[367\]
+ net1018 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_85_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07626_ _03713_ _03730_ net510 vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__mux2_1
XANTENNA__06887__C1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05785__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07557_ net505 net451 _02630_ net443 vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__and4_1
XANTENNA__08628__B1 _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__B net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout620_A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_33_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06508_ net1082 _02612_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_137_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11526__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07488_ net975 _03585_ _03586_ net1068 vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09227_ net569 _04791_ net419 net341 net1600 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__a32o_1
X_06439_ core.register_file.registers_state\[857\] core.register_file.registers_state\[889\]
+ net712 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__mux2_1
XANTENNA__07851__A1 core.decoder.inst\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1150_X net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10309__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07966__X _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09158_ _04924_ net351 net343 net1884 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__a22o_1
X_08109_ net487 _03764_ _03798_ _04209_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__o311a_1
XANTENNA__07064__C1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__A3 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09089_ net2245 net363 net351 _04776_ vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ clknet_leaf_105_clk _00632_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[592\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05614__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05927__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold870 core.register_file.registers_state\[448\] vssd1 vssd1 vccd1 vccd1 net2189
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 core.register_file.registers_state\[102\] vssd1 vssd1 vccd1 vccd1 net2200
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold892 core.register_file.registers_state\[684\] vssd1 vssd1 vccd1 vccd1 net2211
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ clknet_leaf_108_clk _00563_ net1140 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[523\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08022__B _03139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10002_ net1667 net540 net519 _05101_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__a22o_1
XANTENNA__09833__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06017__S1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08867__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10904_ clknet_leaf_4_clk _00416_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[376\]
+ sky130_fd_sc_hd__dfrtp_1
X_11884_ clknet_leaf_53_clk _01353_ net1304 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10835_ clknet_leaf_97_clk _00347_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[307\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05550__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08692__B _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08095__A1 _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10766_ clknet_leaf_89_clk _00278_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[238\]
+ sky130_fd_sc_hd__dfrtp_1
X_10697_ clknet_leaf_40_clk _00209_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[169\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05853__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07055__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05605__B1 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06948__A3 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05837__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06432__S net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ clknet_leaf_61_clk _00830_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[790\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09347__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11249_ clknet_leaf_74_clk _00761_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[721\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09028__B net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06168__A1_N net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05369__C1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05810_ net1060 core.register_file.registers_state\[82\] core.register_file.registers_state\[114\]
+ net690 net648 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__o221a_1
X_06790_ net971 _02893_ _02894_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__or3_1
XANTENNA__06581__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05741_ net1063 core.register_file.registers_state\[180\] net691 core.register_file.registers_state\[148\]
+ net649 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08460_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__inv_2
XANTENNA__05291__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__C1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05672_ net633 _01769_ _01776_ net720 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07411_ core.register_file.registers_state\[536\] core.register_file.registers_state\[568\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08391_ _04482_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11552__RESET_B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07342_ _01664_ _02534_ _02599_ net537 vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08094__S net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10573__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ net996 core.register_file.registers_state\[64\] net890 core.register_file.registers_state\[96\]
+ net829 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_14_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06192__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09012_ net611 _04769_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06224_ net944 core.register_file.registers_state\[581\] net702 core.register_file.registers_state\[613\]
+ net657 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 core.register_file.registers_state\[31\] vssd1 vssd1 vccd1 vccd1 net1419
+ sky130_fd_sc_hd__dlygate4sd3_1
X_06155_ net948 core.register_file.registers_state\[967\] net706 core.register_file.registers_state\[999\]
+ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold111 core.register_file.registers_state\[7\] vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 core.ADR_I\[18\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold133 core.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10196__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold144 core.ADR_I\[28\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05747__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold155 core.ADR_I\[14\] vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
X_06086_ core.register_file.registers_state\[137\] core.register_file.registers_state\[169\]
+ net699 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold166 core.CPU_DAT_I\[18\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold177 _01222_ vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold188 core.CPU_DAT_I\[7\] vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ core.control_logic.instruction\[3\] core.CPU_DAT_O\[3\] net892 vssd1 vssd1
+ vccd1 vccd1 _01067_ sky130_fd_sc_hd__mux2_1
Xfanout602 _04897_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold199 _01205_ vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 net615 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1110_A core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_2
XANTENNA__09889__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 _01521_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1208_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 net650 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ net1122 net601 net383 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__or3b_1
Xfanout657 net659 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_4
XANTENNA__11079__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout668 net680 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout570_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout668_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07995__S1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ _05018_ net293 net259 net1715 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06572__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06988_ core.register_file.registers_state\[265\] core.register_file.registers_state\[297\]
+ core.register_file.registers_state\[393\] core.register_file.registers_state\[425\]
+ net872 net1074 vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux4_1
XANTENNA__05482__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06572__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ core.IO_mod.input_reg\[14\] net253 net728 vssd1 vssd1 vccd1 vccd1 _04788_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05939_ _02040_ _02043_ net629 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08313__A2 _04401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08658_ _04717_ _04728_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__and3_4
XANTENNA__06324__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07521__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07609_ net454 _03319_ net446 net507 vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08589_ core.decoder.inst\[11\] net1117 net742 net611 _04662_ vssd1 vssd1 vccd1 vccd1
+ _04664_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_25_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10620_ clknet_leaf_39_clk _00132_ net1218 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10551_ clknet_leaf_22_clk _00063_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09828__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10482_ net1412 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout992_X net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10187__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06486__S1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ clknet_leaf_15_clk _00615_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[575\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09329__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06260__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08968__A _04860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09563__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07872__A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ clknet_leaf_7_clk _00546_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[506\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08001__A1 _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07591__B _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06563__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05392__A core.decoder.inst\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09501__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07738__S1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05669__A3 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ clknet_leaf_54_clk _01336_ net1300 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10818_ clknet_leaf_78_clk _00330_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[290\]
+ sky130_fd_sc_hd__dfrtp_1
X_11798_ clknet_leaf_31_clk _00009_ net1206 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07276__C1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11630__Q core.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10749_ clknet_leaf_18_clk _00261_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[221\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06951__A _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07766__B net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08240__A1 _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07960_ _03027_ _03402_ _03025_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08878__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06911_ net820 _03012_ _03011_ net785 vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07891_ _01827_ _02747_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__nor2_1
X_09630_ net2475 net393 _05076_ net1001 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__a22o_1
X_06842_ net991 core.register_file.registers_state\[207\] net877 core.register_file.registers_state\[239\]
+ net808 vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a221o_1
XANTENNA__06554__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ net204 net2459 net303 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__mux2_1
X_06773_ net1093 core.register_file.registers_state\[80\] core.register_file.registers_state\[112\]
+ net833 net804 vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__o221a_1
XANTENNA__10939__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08512_ core.pc.current_pc\[26\] _04583_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__nor2_1
X_05724_ net1065 core.register_file.registers_state\[980\] core.register_file.registers_state\[1012\]
+ net692 net1023 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06306__A1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09492_ net603 net204 net316 net261 net2140 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__a32o_1
XANTENNA__10102__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08443_ core.pc.current_pc\[20\] _02779_ net575 vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05655_ net949 core.register_file.registers_state\[694\] net763 vssd1 vssd1 vccd1
+ vccd1 _01760_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ net230 _04466_ _04467_ _04462_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__o31ai_1
XANTENNA__08059__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05586_ net1043 core.register_file.registers_state\[475\] vssd1 vssd1 vccd1 vccd1
+ _01691_ sky130_fd_sc_hd__or2_1
XANTENNA__09256__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07325_ _03426_ _03427_ _03429_ _03428_ net784 net803 vssd1 vssd1 vccd1 vccd1 _03430_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_119_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1060_A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout416_A net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05817__B1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ core.register_file.registers_state\[928\] core.register_file.registers_state\[896\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06861__A _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06207_ net960 _02305_ _02306_ _02311_ net1005 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a311o_1
XANTENNA__10686__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06490__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ net533 _03291_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10169__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06138_ net1054 core.register_file.registers_state\[135\] vssd1 vssd1 vccd1 vccd1
+ _02243_ sky130_fd_sc_hd__or2_1
XANTENNA__07034__A2 _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08782__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06069_ _02154_ _02160_ _02173_ net721 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_4
XANTENNA_fanout1113_X net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06793__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_4
Xfanout432 net435 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
Xfanout443 net447 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_2
XANTENNA__07417__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout952_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout465 _04709_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_4
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout487 net488 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
X_09828_ net219 net2171 net380 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_2
X_09759_ _04987_ net286 net257 net1555 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09495__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11403__RESET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08954__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11721_ clknet_leaf_36_clk _01233_ net1219 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11652_ clknet_leaf_36_clk _01164_ net1219 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09247__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07258__C1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10603_ clknet_leaf_110_clk _00115_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09798__A1 _04812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11583_ clknet_leaf_27_clk _01095_ net1204 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05808__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09558__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10534_ clknet_leaf_100_clk _00046_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06771__A _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11244__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05284__B2 _01395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06481__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07586__B _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10465_ net1411 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08034__Y _04139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07078__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10396_ net1322 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07576__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11017_ clknet_leaf_39_clk _00529_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[489\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09486__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11144__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_0_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07497__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05440_ net1048 core.register_file.registers_state\[478\] core.register_file.registers_state\[510\]
+ net674 net1014 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06157__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09238__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05371_ core.register_file.registers_state\[798\] core.register_file.registers_state\[830\]
+ core.register_file.registers_state\[926\] core.register_file.registers_state\[958\]
+ net881 net1075 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07110_ net1086 _03213_ _03214_ net1068 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08090_ _03716_ _03726_ net486 vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload20 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_8
X_07041_ _03052_ _03055_ _03083_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload31 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__inv_8
Xclkload42 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload53 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__clkinv_8
Xclkload64 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_45_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11737__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload75 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__clkinv_2
Xclkload86 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload97 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_6
XANTENNA__06224__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07421__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10020__B2 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08992_ net744 net465 _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__and3_1
X_07943_ _03658_ _03820_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nor2_1
XANTENNA__10761__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ _03713_ _03774_ _03976_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_108_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09931__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ _04982_ net395 net391 net1832 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__a22o_1
X_06825_ _02921_ _02922_ _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09544_ _04889_ core.register_file.registers_state\[586\] net303 vssd1 vssd1 vccd1
+ vccd1 _00626_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09477__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06756_ net781 _02853_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_65_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07451__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05707_ net1056 core.register_file.registers_state\[53\] net756 vssd1 vssd1 vccd1
+ vccd1 _01812_ sky130_fd_sc_hd__and3_1
X_09475_ _04981_ net315 net261 net1781 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a22o_1
X_06687_ net1099 core.register_file.registers_state\[723\] core.register_file.registers_state\[755\]
+ net840 net817 vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout533_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09492__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ _04496_ _04513_ _04512_ _04505_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__o211a_2
XFILLER_0_47_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09229__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05638_ _01741_ _01742_ net1026 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11267__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ _02085_ _04450_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05569_ net937 core.register_file.registers_state\[827\] net758 net922 vssd1 vssd1
+ vccd1 vccd1 _01674_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout1063_X net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__inv_6
XFILLER_0_89_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07308_ _02905_ _03412_ _02786_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07687__A _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08452__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08288_ _04376_ _04379_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05478__Y _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07239_ net1107 core.register_file.registers_state\[129\] net847 core.register_file.registers_state\[161\]
+ net826 vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__o221a_1
XANTENNA__10317__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10250_ net1126 net1435 net910 _05233_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06215__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07693__Y _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A1 core.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__B1_N _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10181_ net108 net917 net907 net1590 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1205 net1207 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1216 net1224 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1227 net1229 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
Xfanout240 _05247_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_4
XFILLER_0_100_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1238 net1239 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05974__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
Xfanout1249 net1250 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout262 _05059_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_4
Xfanout273 _05086_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_4
XANTENNA__08063__S0 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout284 _05081_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_6
Xfanout295 net298 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09841__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09180__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07191__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08965__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09468__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07214__X _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ clknet_leaf_72_clk _01216_ net1271 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08691__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11635_ clknet_leaf_71_clk _01147_ net1270 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09288__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ clknet_leaf_26_clk _01078_ net1203 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10250__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06454__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10517_ clknet_leaf_36_clk _00029_ net1221 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11497_ clknet_leaf_38_clk _01009_ net1213 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[969\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08205__B _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10448_ net1427 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10784__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__B2 _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10379_ net1343 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09036__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06509__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__B1 _03810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05980__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06509__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__C1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06610_ _02713_ _02714_ net1089 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07590_ _02384_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_103_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09459__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06390__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10069__A1 _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06541_ net772 _02640_ _02645_ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ net2448 net207 net337 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06472_ net1034 core.register_file.registers_state\[728\] core.register_file.registers_state\[760\]
+ net665 net651 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08891__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ _03685_ _04187_ _04309_ _04315_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05496__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05423_ net1048 core.register_file.registers_state\[862\] core.register_file.registers_state\[894\]
+ net678 net1027 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05496__B2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09191_ _04987_ net351 net423 net1601 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08142_ _03390_ _03391_ _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__o21ai_1
X_05354_ _01388_ _01390_ _01393_ _01395_ net1070 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__o221a_4
XANTENNA__09631__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08073_ _02345_ _03231_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05285_ core.decoder.inst\[12\] _01397_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08115__B _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06996__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06996__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07024_ net807 _03127_ _03128_ net1084 vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a211o_1
XANTENNA__09926__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05458__C net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09934__A1 core.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06748__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1023_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08975_ net566 _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout483_A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 core.register_file.registers_state\[933\] vssd1 vssd1 vccd1 vccd1 net1334
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 core.register_file.registers_state\[1009\] vssd1 vssd1 vccd1 vccd1 net1345
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 core.register_file.registers_state\[951\] vssd1 vssd1 vccd1 vccd1 net1356
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _01987_ _02873_ net548 _01958_ net900 vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__a32o_1
XANTENNA__09698__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold48 core.SEL_I\[0\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 core.register_file.registers_state\[1006\] vssd1 vssd1 vccd1 vccd1 net1378
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09162__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ net532 _03959_ _03961_ _03657_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout650_A _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__B net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ core.register_file.registers_state\[781\] core.register_file.registers_state\[813\]
+ net865 vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__mux2_1
XANTENNA__05723__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07788_ net497 _03675_ _03799_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06586__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07034__X _03139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ _04857_ net396 net307 net1761 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a22o_1
X_06739_ _01926_ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout915_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1278_X net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09458_ _04950_ net316 net311 net2015 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a22o_1
XANTENNA__09870__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08409_ _04498_ _04499_ net598 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09389_ net2109 net327 net316 _04839_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11420_ clknet_leaf_42_clk _00932_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08976__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ clknet_leaf_8_clk _00863_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06987__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06531__S0 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10302_ net26 net902 net796 net2470 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_56_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09836__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11282_ clknet_leaf_68_clk _00794_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[754\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08728__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ net77 net915 vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10164_ net1125 net1367 net910 _05206_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__a31o_1
XANTENNA_input44_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 _01368_ vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_4
XANTENNA__08679__C _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06203__A3 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1013 net1016 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_4
Xfanout1024 core.decoder.inst\[22\] vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_37_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05384__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1046 net1050 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
X_10095_ _04043_ net557 net590 core.pc.current_pc\[17\] net472 vssd1 vssd1 vccd1 vccd1
+ _05157_ sky130_fd_sc_hd__o221a_1
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09689__A0 _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1068 core.decoder.inst\[18\] vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1081 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06199__C net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09153__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11432__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06911__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ clknet_leaf_62_clk _00509_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[469\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07011__S1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06124__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05478__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11618_ clknet_leaf_31_clk _01130_ net1205 vssd1 vssd1 vccd1 vccd1 core.READ_I sky130_fd_sc_hd__dfrtp_2
XFILLER_0_113_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__A _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08967__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11549_ clknet_leaf_18_clk _01061_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1021\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold507 core.register_file.registers_state\[268\] vssd1 vssd1 vccd1 vccd1 net1826
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__S net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold518 core.register_file.registers_state\[235\] vssd1 vssd1 vccd1 vccd1 net1837
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 core.register_file.registers_state\[348\] vssd1 vssd1 vccd1 vccd1 net1848
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08195__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05294__B core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 core.register_file.registers_state\[471\] vssd1 vssd1 vccd1 vccd1 net2526
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ net606 net215 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__and2_1
Xhold1218 wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
X_05972_ net1036 core.register_file.registers_state\[973\] core.register_file.registers_state\[1005\]
+ net665 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1229 core.register_file.registers_state\[699\] vssd1 vssd1 vccd1 vccd1 net2548
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08886__A core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ _03451_ _03478_ _03814_ net527 vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08691_ net730 _04140_ _04755_ net525 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a211o_2
XANTENNA__07155__B2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07642_ net452 _03023_ net444 net501 vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07573_ _03673_ _03676_ net482 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09312_ _04935_ net421 net333 net2141 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__a22o_1
X_06524_ _02619_ _02622_ _02628_ net968 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06115__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07458__A2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09852__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05469__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05469__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ net558 _04846_ _05037_ net339 net2058 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__a32o_1
X_06455_ net723 _02546_ _02558_ _02559_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a22o_4
XFILLER_0_106_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06761__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_A _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05406_ core.decoder.inst\[24\] net749 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__and2_4
XFILLER_0_12_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09174_ _04956_ net352 net343 net2128 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__a22o_1
X_06386_ _02489_ _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__and2_1
XANTENNA__08126__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10214__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05337_ net1315 net1911 _01442_ core.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 _00005_
+ sky130_fd_sc_hd__a22o_1
X_08125_ _03898_ _04131_ net531 vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1140_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06513__S0 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07091__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05268_ core.pc.current_pc\[23\] vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
X_08056_ _04138_ _04160_ net478 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05641__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout698_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ net539 _02524_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09907__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09383__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05929__C1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08591__B1 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ net2393 net367 _04945_ net432 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07909_ net486 _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ net2540 net370 _04899_ net439 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10330__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ clknet_leaf_12_clk _00432_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[392\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05280__A_N core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05424__S net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ clknet_leaf_73_clk _00363_ net1272 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[323\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09843__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ clknet_leaf_97_clk _00294_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[254\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06255__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08949__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ clknet_leaf_110_clk _00915_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[875\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05880__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09071__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ clknet_leaf_99_clk _00846_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07621__A2 _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11265_ clknet_leaf_86_clk _00777_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[737\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05395__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ net1127 net1448 net912 _05216_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a31o_1
XANTENNA__08031__C1 _04135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08177__A3 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ clknet_leaf_41_clk _00708_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[668\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07385__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07385__B2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ core.pc.current_pc\[30\] _05187_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10078_ core.pc.current_pc\[11\] net590 vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__or2_1
XANTENNA__07137__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10141__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05699__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10972__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A0 _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08637__A1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09330__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_06240_ net583 _02343_ _02344_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a21o_2
XFILLER_0_26_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05871__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05289__B core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06171_ net554 _02273_ _02275_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05871__B2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09601__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold304 core.register_file.registers_state\[272\] vssd1 vssd1 vccd1 vccd1 net1623
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold315 core.register_file.registers_state\[778\] vssd1 vssd1 vccd1 vccd1 net1634
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 core.register_file.registers_state\[392\] vssd1 vssd1 vccd1 vccd1 net1645
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold337 core.register_file.registers_state\[780\] vssd1 vssd1 vccd1 vccd1 net1656
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold348 core.CPU_DAT_I\[11\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05623__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09930_ core.decoder.inst\[19\] core.CPU_DAT_O\[19\] net892 vssd1 vssd1 vccd1 vccd1
+ _01083_ sky130_fd_sc_hd__mux2_1
Xhold359 core.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 net807 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09861_ _04929_ net387 net267 net2084 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__a22o_1
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout828 net830 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_4
Xfanout839 net846 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload16_A clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ net727 _03839_ net525 _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a211o_1
X_09792_ _04782_ net385 net273 net1725 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__a22o_1
Xhold1004 core.register_file.registers_state\[127\] vssd1 vssd1 vccd1 vccd1 net2323
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 core.register_file.registers_state\[863\] vssd1 vssd1 vccd1 vccd1 net2334
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 core.register_file.registers_state\[339\] vssd1 vssd1 vccd1 vccd1 net2345
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08743_ net564 net606 net218 vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and3_1
Xhold1037 core.register_file.registers_state\[121\] vssd1 vssd1 vccd1 vccd1 net2356
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 core.register_file.registers_state\[64\] vssd1 vssd1 vccd1 vccd1 net2367
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05955_ net616 _02054_ _02056_ net631 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a31o_1
Xhold1059 core.register_file.registers_state\[185\] vssd1 vssd1 vccd1 vccd1 net2378
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09999__X _05100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__A2 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ net2097 net467 net433 _04743_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__a22o_1
XANTENNA__10003__X _05102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06336__C1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05886_ net963 _01990_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _03721_ _03729_ net493 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout446_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05785__S1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07556_ _01488_ net498 net451 net443 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__and4b_1
XANTENNA__08628__A1 core.IO_mod.input_reg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06507_ core.register_file.registers_state\[285\] core.register_file.registers_state\[317\]
+ core.register_file.registers_state\[413\] core.register_file.registers_state\[445\]
+ net868 net1070 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07487_ net972 _03590_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout613_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09226_ _04787_ net416 net339 net1734 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06438_ core.register_file.registers_state\[985\] core.register_file.registers_state\[1017\]
+ net712 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__mux2_1
XANTENNA__07851__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ _04922_ net354 net344 net2082 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06369_ net1059 core.register_file.registers_state\[642\] vssd1 vssd1 vccd1 vccd1
+ _02474_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08108_ net491 _04161_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__a21o_1
XANTENNA__07064__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ net2210 net363 net353 _04770_ vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout982_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05614__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08039_ net532 _04016_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__nor2_1
XANTENNA__10325__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold860 core.register_file.registers_state\[635\] vssd1 vssd1 vccd1 vccd1 net2179
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 core.register_file.registers_state\[486\] vssd1 vssd1 vccd1 vccd1 net2190
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11081__RESET_B net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold882 core.register_file.registers_state\[469\] vssd1 vssd1 vccd1 vccd1 net2201
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08159__A3 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold893 core.register_file.registers_state\[374\] vssd1 vssd1 vccd1 vccd1 net2212
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ clknet_leaf_1_clk _00562_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[522\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06104__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ net724 _02145_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__and2_2
XANTENNA__09108__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06327__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06878__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10903_ clknet_leaf_22_clk _00415_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[375\]
+ sky130_fd_sc_hd__dfrtp_1
X_11883_ clknet_leaf_48_clk _01352_ net1312 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09816__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10834_ clknet_leaf_69_clk _00346_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[306\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08465__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10765_ clknet_leaf_0_clk _00277_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[237\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10696_ clknet_leaf_95_clk _00208_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05853__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09044__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09595__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05605__A1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11317_ clknet_leaf_63_clk _00829_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06948__A4 _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08213__B _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ clknet_leaf_105_clk _00760_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[720\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08555__B1 _01508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09898__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap411_A _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ clknet_leaf_108_clk _00691_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[651\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06566__C1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05740_ _01843_ _01844_ net718 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05671_ net965 _01770_ _01775_ net629 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a211o_1
X_07410_ core.register_file.registers_state\[600\] core.register_file.registers_state\[632\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11150__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08390_ _01988_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__or2_1
XANTENNA__05541__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09060__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ _03433_ _03445_ net771 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__mux2_8
XFILLER_0_9_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09283__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06097__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07272_ net814 _03375_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09011_ net2040 net428 _04980_ net434 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__a22o_1
XANTENNA__05844__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06192__S1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06223_ net1029 _02324_ _02327_ net633 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__o211a_1
XANTENNA__09035__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07046__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06154_ net633 _02258_ net723 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08243__C1 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold101 core.register_file.registers_state\[1001\] vssd1 vssd1 vccd1 vccd1 net1420
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09586__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06623__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold112 core.register_file.registers_state\[15\] vssd1 vssd1 vccd1 vccd1 net1431
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 core.ADR_I\[11\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 core.IO_mod.data_from_mem\[30\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06085_ _02185_ _02189_ net1005 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a21oi_1
Xhold145 net161 vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 net185 vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold167 _01219_ vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09934__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ core.control_logic.instruction\[2\] core.CPU_DAT_O\[2\] net892 vssd1 vssd1
+ vccd1 vccd1 _01066_ sky130_fd_sc_hd__mux2_1
Xhold178 core.register_file.registers_state\[1019\] vssd1 vssd1 vccd1 vccd1 net1497
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold189 _01208_ vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _04706_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07349__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 net637 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_4
Xfanout647 net650 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_4
X_09844_ net242 net2334 net381 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_2
XANTENNA__10353__A0 _05105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1103_A core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout669 net680 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07307__X _03412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ net603 net203 net288 net257 net1586 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__a32o_1
X_06987_ net791 _03088_ _03091_ net775 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout563_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08726_ net1834 net466 net431 _04787_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__a22o_1
X_05938_ net625 _02041_ _02042_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_83_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ net729 _04200_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout730_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05869_ _01972_ _01973_ net623 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout828_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1093_X net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07608_ _03705_ _03712_ net496 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08588_ net746 net611 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07539_ net480 _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nor2_1
XANTENNA__07809__C1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09274__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10550_ clknet_leaf_59_clk _00062_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07202__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09209_ _05020_ net356 net424 net1644 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__a22o_1
XANTENNA__05835__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10481_ net1432 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09026__B2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08234__C1 _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09577__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05938__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06260__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ clknet_leaf_93_clk _00614_ net1239 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[574\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09844__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09329__A2 _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold690 core.register_file.registers_state\[873\] vssd1 vssd1 vccd1 vccd1 net2009
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11023__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08968__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11033_ clknet_leaf_55_clk _00545_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[505\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10344__A0 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__C1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06769__A _01987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09501__A2 _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11866_ clknet_leaf_52_clk _01335_ net1302 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06720__C1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10817_ clknet_leaf_83_clk _00329_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[289\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11797_ clknet_leaf_31_clk _00008_ net1201 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08208__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06079__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09804__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06079__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10748_ clknet_leaf_39_clk _00260_ net1218 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05826__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05826__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09017__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10679_ clknet_leaf_21_clk _00191_ net1182 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[151\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09568__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09039__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08240__A2 _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08878__B _04860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06910_ _03013_ _03014_ net790 vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__o21a_1
XANTENNA__10335__A0 _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07890_ _03774_ _03856_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nor2_1
XANTENNA__06679__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__Y _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07200__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ net991 core.register_file.registers_state\[79\] net877 core.register_file.registers_state\[111\]
+ net826 vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _04893_ net2374 net303 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06772_ core.register_file.registers_state\[16\] core.register_file.registers_state\[48\]
+ core.register_file.registers_state\[144\] core.register_file.registers_state\[176\]
+ net865 net817 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_121_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05762__B1 core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08894__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ core.pc.current_pc\[26\] _04583_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__and2_1
X_05723_ net1052 net899 _01507_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a21oi_2
X_09491_ _05012_ net316 net261 net1876 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a22o_1
XANTENNA__11666__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08700__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08442_ core.pc.current_pc\[19\] _04529_ net600 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05654_ net1056 net753 core.register_file.registers_state\[662\] vssd1 vssd1 vccd1
+ vccd1 _01759_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07303__A _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08373_ _04464_ _04465_ _04451_ _04455_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08059__A2 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09256__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05585_ net939 core.register_file.registers_state\[507\] net759 vssd1 vssd1 vccd1
+ vccd1 _01690_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07797__X _03902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09929__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ core.register_file.registers_state\[91\] core.register_file.registers_state\[123\]
+ net866 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__mux2_1
XANTENNA__10690__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07255_ net1089 _03355_ _03356_ _03359_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout311_A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09008__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_A core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05758__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06206_ net1013 _02308_ _02310_ net1027 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__o211a_1
XANTENNA__07449__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07186_ net504 net492 net477 _01632_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a31o_1
X_06137_ _02206_ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1220_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06778__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06242__A1 core.decoder.inst\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06242__B2 core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06068_ _02164_ _02167_ _02169_ _02172_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout680_A _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 net402 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_4
XANTENNA__07990__A1 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05450__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_A _01463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _05029_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07692__B _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10326__A0 _05111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 net435 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_4
Xfanout444 net446 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_2
XANTENNA__07417__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 _02529_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1106_X net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09192__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 _04667_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_8
Xfanout477 net481 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ net220 net2268 net380 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
XANTENNA__09731__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_2
Xfanout499 net503 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout945_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07742__B2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ _04985_ net291 net260 net1656 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__a22o_1
XANTENNA__05753__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08709_ core.IO_mod.data_from_mem\[11\] net248 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _04888_ net2389 net278 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__mux2_1
X_11720_ clknet_leaf_54_clk net1482 net1299 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05505__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ clknet_leaf_54_clk _01163_ net1300 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09247__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07258__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ clknet_leaf_111_clk _00114_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09839__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09798__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11582_ clknet_leaf_27_clk _01094_ net1204 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10533_ clknet_leaf_92_clk _00045_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05668__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ net1396 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08222__A2 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10395_ net1447 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07430__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07981__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05674__Y _01779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10317__A0 _05102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08050__Y _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06499__A _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09183__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ clknet_leaf_14_clk _00528_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[488\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09722__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07733__A1 _03697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05744__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10096__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06438__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08219__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ clknet_leaf_24_clk net44 net1183 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05370_ _01467_ net772 _01474_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__or3_2
XANTENNA__09789__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11069__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinvlp_4
X_07040_ _03115_ _03144_ _03087_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__and3b_1
Xclkload21 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__06472__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload32 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__inv_8
XANTENNA__06472__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload43 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_8
Xclkload54 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload65 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__inv_6
XFILLER_0_80_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload76 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__inv_8
Xclkload87 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_12
XANTENNA__09410__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload98 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__inv_16
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06224__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10020__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06901__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ net614 net224 vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07942_ _03056_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__xor2_2
XFILLER_0_103_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10308__A0 _02421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07873_ _01746_ net552 _03618_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__a211o_1
XANTENNA__06202__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07724__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ _04980_ net398 net392 net1935 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06824_ net779 _02925_ _02928_ net767 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_69_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06932__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09543_ _04888_ net2426 net306 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06755_ net778 _02856_ _02859_ net773 vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_65_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout359_A net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05706_ _01807_ _01810_ net629 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07488__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _04979_ net319 net262 net2008 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a22o_1
X_06686_ net1099 core.register_file.registers_state\[595\] core.register_file.registers_state\[627\]
+ net840 net805 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08425_ _04496_ _04513_ _04505_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o21a_1
X_05637_ net1040 core.register_file.registers_state\[471\] core.register_file.registers_state\[503\]
+ net671 net1010 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1170_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1268_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08356_ _02085_ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05568_ net937 core.register_file.registers_state\[955\] net757 net1012 vssd1 vssd1
+ vccd1 vccd1 _01673_ sky130_fd_sc_hd__o31a_1
XFILLER_0_80_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload4 clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_8
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07307_ _03403_ _03407_ _03411_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__a21o_2
XANTENNA__07687__B _01550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ _04386_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05499_ core.register_file.registers_state\[540\] core.register_file.registers_state\[572\]
+ net707 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1056_X net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06463__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07179__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07238_ core.register_file.registers_state\[33\] core.register_file.registers_state\[1\]
+ net847 vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05671__C1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09401__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07169_ _03272_ _03273_ net976 vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07907__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10180_ net1651 net916 net906 net1648 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a22o_1
XANTENNA__10586__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05423__C1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1207 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10333__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1217 net1224 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_4
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
Xfanout241 _04880_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07990__X _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09165__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1239 net1250 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__buf_2
XANTENNA__05427__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout274 _05083_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_8
Xfanout285 _05081_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_2
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net298 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_4
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06923__C1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ clknet_leaf_70_clk net2496 net1275 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11211__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11634_ clknet_leaf_52_clk _01146_ net1302 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06782__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11565_ clknet_leaf_33_clk _01077_ net1205 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07597__B _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05398__A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06454__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10516_ clknet_leaf_36_clk _00028_ net1221 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11361__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11496_ clknet_leaf_9_clk _01008_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[968\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_126_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10447_ net1414 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06206__A1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10378_ net1366 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__05414__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09156__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06914__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06390__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10069__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06540_ net1087 _02641_ _02644_ net780 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06471_ net1034 core.register_file.registers_state\[984\] core.register_file.registers_state\[1016\]
+ net665 net1008 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__o221a_1
XANTENNA__06142__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08682__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _03819_ _03980_ _04310_ _04312_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06693__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05422_ net627 _01525_ _01526_ net720 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_116_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09190_ _04985_ net354 net424 net1826 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__a22o_1
XANTENNA__05800__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ _03390_ _03391_ net528 vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05353_ _01387_ _01389_ _01392_ _01394_ net987 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a221o_2
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06445__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ net1112 _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05284_ _01388_ _01390_ _01393_ _01395_ core.decoder.inst\[12\] vssd1 vssd1 vccd1
+ vccd1 _01399_ sky130_fd_sc_hd__o221a_4
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07023_ net988 core.register_file.registers_state\[680\] net872 core.register_file.registers_state\[648\]
+ net821 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__o221a_1
XFILLER_0_109_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08198__A1 _03788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09395__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11521__SET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ _04870_ net601 vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1016_A core.decoder.inst\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09147__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 core.register_file.registers_state\[963\] vssd1 vssd1 vccd1 vccd1 net1335
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _02902_ _02906_ _03410_ net528 vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a31oi_1
Xhold27 core.register_file.registers_state\[928\] vssd1 vssd1 vccd1 vccd1 net1346
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 core.register_file.registers_state\[998\] vssd1 vssd1 vccd1 vccd1 net1357
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 core.register_file.registers_state\[959\] vssd1 vssd1 vccd1 vccd1 net1368
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ net487 _03910_ _03960_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__a21o_1
XANTENNA__05708__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06807_ core.register_file.registers_state\[909\] core.register_file.registers_state\[941\]
+ net863 vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__mux2_1
X_07787_ net497 _03675_ _03799_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout643_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09526_ _04851_ net401 net310 net1976 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06738_ _01957_ _01987_ _02526_ _02527_ net538 vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__o41a_1
XFILLER_0_52_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07969__Y _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09457_ _04948_ net325 net314 net2241 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a22o_1
X_06669_ net1109 core.register_file.registers_state\[468\] core.register_file.registers_state\[500\]
+ net859 net1080 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout810_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06133__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07330__C1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08408_ core.pc.current_pc\[15\] _04477_ core.pc.current_pc\[16\] vssd1 vssd1 vccd1
+ vccd1 _04499_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06684__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06684__B2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ net2029 net329 net322 _04833_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08339_ _04433_ _04434_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10328__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11350_ clknet_leaf_61_clk _00862_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08830__C1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05649__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ net25 net905 _05244_ core.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 _01298_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06531__S1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05644__C1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ clknet_leaf_73_clk _00793_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[753\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09386__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ net1128 net1425 net913 _05224_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10163_ net136 net914 vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__and2_1
Xfanout1003 _01365_ vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1014 net1016 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__buf_2
Xfanout1025 net1033 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__buf_4
Xfanout1036 net1038 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input37_A gpio_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1050 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
X_10094_ net473 _05155_ _05156_ net517 net1625 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__a32o_1
Xfanout1058 core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_4
Xfanout1069 net1072 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_4
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06372__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10601__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ clknet_leaf_51_clk _00508_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05580__D1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08992__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09310__B1 _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07879__Y _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05478__A2 _01582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11617_ clknet_leaf_33_clk _01129_ net1205 vssd1 vssd1 vccd1 vccd1 core.i_hit sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10758__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08216__B _04317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11548_ clknet_leaf_43_clk _01060_ net1283 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1020\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_53_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold508 core.register_file.registers_state\[47\] vssd1 vssd1 vccd1 vccd1 net1827
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold519 core.register_file.registers_state\[710\] vssd1 vssd1 vccd1 vccd1 net1838
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11479_ clknet_leaf_6_clk _00991_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[951\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11107__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09377__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09129__A0 _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06060__C1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1208 core.register_file.registers_state\[202\] vssd1 vssd1 vccd1 vccd1 net2527
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05971_ net1036 core.register_file.registers_state\[845\] core.register_file.registers_state\[877\]
+ net665 net923 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__o221a_1
XANTENNA__11257__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1219 core.register_file.registers_state\[313\] vssd1 vssd1 vccd1 vccd1 net2538
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08886__B net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07710_ _03478_ _03814_ _03451_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_105_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08690_ _04701_ _04717_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07641_ _03744_ _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07572_ _03676_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09311_ net561 _04933_ _05048_ net334 net2546 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a32o_1
XANTENNA__09301__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06523_ net970 _02626_ _02627_ _02625_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__o31a_1
XFILLER_0_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09242_ core.register_file.registers_state\[312\] net474 net544 vssd1 vssd1 vccd1
+ vccd1 _05037_ sky130_fd_sc_hd__o21a_1
XANTENNA__06666__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06454_ net635 _02552_ _02553_ net719 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__o31a_1
XFILLER_0_8_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05405_ net896 _01408_ _01410_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06761__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09173_ _04954_ net355 net344 net2096 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06385_ net944 core.register_file.registers_state\[961\] net702 core.register_file.registers_state\[993\]
+ net927 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout224_A _04730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09937__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ _04022_ _04041_ _04223_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__o211a_4
XANTENNA__06418__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05336_ net1315 net1691 core.ru.state\[4\] _01442_ vssd1 vssd1 vccd1 vccd1 _00004_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08841__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09080__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05626__C1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06513__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _03722_ _03723_ net500 vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux2_1
XANTENNA__07091__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05267_ core.pc.current_pc\[19\] vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1133_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ net768 _03110_ _03098_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__o21a_4
XANTENNA__09368__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05641__A2 _01745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout593_A _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A1 _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07379__C1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A0 _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1300_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout760_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ net565 _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout858_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _03634_ _03642_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ net573 net207 net737 vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_32_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07839_ net529 _03918_ _03919_ _03941_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a31o_1
XANTENNA__06354__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ clknet_leaf_78_clk _00362_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[322\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09509_ _04760_ net398 net308 net1777 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__a22o_1
X_10781_ clknet_leaf_17_clk _00293_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[253\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05865__C1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10851__RESET_B net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06409__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11402_ clknet_leaf_1_clk _00914_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[874\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09071__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11333_ clknet_leaf_87_clk _00845_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07875__B _03697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09359__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11264_ clknet_leaf_59_clk _00776_ net1286 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[736\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08052__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10215_ net99 net915 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__and2_1
X_11195_ clknet_leaf_21_clk _00707_ net1190 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06188__A3 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__A _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _05193_ _05194_ net556 vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10077_ net1509 net517 _05145_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__a21o_1
XANTENNA__09531__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10141__A1 _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06345__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06440__S0 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10979_ clknet_leaf_71_clk _00491_ net1270 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[451\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06648__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06648__B2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__B net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06112__A3 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09598__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06170_ net585 _02274_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07785__B _03763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 core.register_file.registers_state\[394\] vssd1 vssd1 vccd1 vccd1 net1624
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold316 core.register_file.registers_state\[280\] vssd1 vssd1 vccd1 vccd1 net1635
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold327 core.register_file.registers_state\[819\] vssd1 vssd1 vccd1 vccd1 net1646
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05586__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 core.register_file.registers_state\[544\] vssd1 vssd1 vccd1 vccd1 net1657
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold349 _01212_ vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06820__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout807 _01460_ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
X_09860_ _04927_ net387 net267 net2183 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__a22o_1
XANTENNA__08897__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net823 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_4
Xfanout829 net830 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08573__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06179__A3 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05873__X _01978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ net726 _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__nor2_1
XANTENNA__09770__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ net563 _04776_ net383 net270 net1947 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__a32o_1
XFILLER_0_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1005 core.register_file.registers_state\[353\] vssd1 vssd1 vccd1 vccd1 net2324
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 core.register_file.registers_state\[669\] vssd1 vssd1 vccd1 vccd1 net2335
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 core.register_file.registers_state\[105\] vssd1 vssd1 vccd1 vccd1 net2346
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11380__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08742_ net606 net218 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__and2_1
X_05954_ _02057_ _02058_ net620 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__o21a_1
Xhold1038 core.register_file.registers_state\[583\] vssd1 vssd1 vccd1 vccd1 net2357
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 core.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09522__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08673_ net568 _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__and2_1
XANTENNA__06336__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05885_ core.register_file.registers_state\[303\] core.register_file.registers_state\[271\]
+ core.register_file.registers_state\[431\] core.register_file.registers_state\[399\]
+ net681 net1018 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_124_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07624_ _03724_ _03728_ net483 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06887__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07555_ net499 _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__or2_2
XFILLER_0_53_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08628__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout341_A _05031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1083_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout439_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ net789 _02607_ _02610_ net776 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__o211a_1
XANTENNA__06639__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07486_ net1100 core.register_file.registers_state\[607\] core.register_file.registers_state\[639\]
+ net844 net806 vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_98_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05847__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ _04782_ net419 net340 net1707 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06437_ core.register_file.registers_state\[793\] core.register_file.registers_state\[825\]
+ net712 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1250_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09589__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09156_ _04920_ net351 net343 net1837 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06368_ net952 core.register_file.registers_state\[706\] net710 core.register_file.registers_state\[738\]
+ net646 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_20_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08107_ _03664_ _04210_ _04211_ _02518_ _03688_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05319_ net1070 net1082 core.decoder.inst\[19\] net1066 vssd1 vssd1 vccd1 vccd1 _01433_
+ sky130_fd_sc_hd__or4_1
XANTENNA__07064__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ net2214 net364 net355 _04764_ vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_110_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06299_ net1062 core.register_file.registers_state\[547\] net754 vssd1 vssd1 vccd1
+ vccd1 _02404_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1136_X net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08038_ _03396_ _04141_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold850 core.register_file.registers_state\[593\] vssd1 vssd1 vccd1 vccd1 net2169
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_A _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 core.register_file.registers_state\[681\] vssd1 vssd1 vccd1 vccd1 net2180
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold872 core.register_file.registers_state\[747\] vssd1 vssd1 vccd1 vccd1 net2191
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 core.register_file.registers_state\[630\] vssd1 vssd1 vccd1 vccd1 net2202
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold894 core.register_file.registers_state\[124\] vssd1 vssd1 vccd1 vccd1 net2213
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11572__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06024__C1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ core.CPU_DAT_I\[10\] net541 net520 _05100_ vssd1 vssd1 vccd1 vccd1 _01142_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09761__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09989_ net1540 net540 net519 _02485_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10341__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06327__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ clknet_leaf_43_clk _00414_ net1286 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[374\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11882_ clknet_leaf_50_clk _01351_ net1307 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ clknet_leaf_75_clk _00345_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[305\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05550__A1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10764_ clknet_leaf_101_clk _00276_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[236\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05838__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10695_ clknet_leaf_91_clk _00207_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05853__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06790__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09044__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_101_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05605__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06802__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11316_ clknet_leaf_56_clk _00828_ net1294 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[788\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06802__B2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08004__B1 _04108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ clknet_leaf_82_clk _00759_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[719\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09752__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09606__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ clknet_leaf_2_clk _00690_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[650\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05369__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ net470 _05177_ _05180_ net515 net1478 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09504__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06030__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06869__A1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05670_ _01772_ _01774_ net1032 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09807__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11488__SET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07340_ net968 _03436_ _03439_ _03441_ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07271_ net1109 core.register_file.registers_state\[128\] net859 core.register_file.registers_state\[160\]
+ net828 vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__o221a_1
XANTENNA__09995__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09010_ net567 net604 _04888_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_132_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06222_ _02325_ _02326_ net963 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08617__A_N _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09035__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06153_ net963 _02256_ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold102 core.register_file.registers_state\[17\] vssd1 vssd1 vccd1 vccd1 net1421
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 core.register_file.registers_state\[1007\] vssd1 vssd1 vccd1 vccd1 net1432
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold124 core.ADR_I\[12\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold135 core.ADR_I\[20\] vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06084_ net641 _02186_ _02188_ net1028 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a211o_1
XANTENNA__11819__Q net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 core.CPU_DAT_I\[12\] vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 core.CPU_DAT_I\[8\] vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold168 core.register_file.registers_state\[1005\] vssd1 vssd1 vccd1 vccd1 net1487
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold179 core.ADR_I\[0\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ core.control_logic.instruction\[1\] core.CPU_DAT_O\[1\] net891 vssd1 vssd1
+ vccd1 vccd1 _01065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout604 _04706_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_2
Xfanout615 _04658_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
Xfanout626 _01523_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_4
XANTENNA__09743__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout637 net642 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_4
X_09843_ net243 net2375 net381 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
Xfanout648 net650 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_4
Xfanout659 net664 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XANTENNA_fanout291_A _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ net785 _03089_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__or3_1
X_09774_ _05015_ net292 net259 net1713 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09950__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05937_ net946 core.register_file.registers_state\[206\] net704 core.register_file.registers_state\[238\]
+ net643 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a221o_1
X_08725_ net564 _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout556_A net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1298_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ core.IO_mod.data_from_mem\[3\] net249 _04727_ vssd1 vssd1 vccd1 vccd1 _04728_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08566__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05868_ net1062 core.register_file.registers_state\[593\] core.register_file.registers_state\[625\]
+ net687 net646 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_54_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ _03708_ _03711_ net485 vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08587_ core.decoder.inst\[11\] net895 _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout723_A _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05799_ net648 _01903_ _01902_ net966 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout1086_X net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07538_ net508 _03640_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06086__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07469_ _03570_ _03573_ net632 vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1253_X net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_69_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09208_ _05018_ net362 net424 net1681 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ net1378 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10812__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09026__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ net210 net2376 net348 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10336__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__B _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10041__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05599__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ clknet_leaf_16_clk _00613_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[573\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold680 core.register_file.registers_state\[314\] vssd1 vssd1 vccd1 vccd1 net1999
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07645__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold691 core.register_file.registers_state\[416\] vssd1 vssd1 vccd1 vccd1 net2010
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ clknet_leaf_5_clk _00544_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[504\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09734__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06548__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__A3 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11468__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06181__D1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11865_ clknet_leaf_54_clk _01334_ net1300 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11841__D net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10816_ clknet_leaf_55_clk _00328_ net1301 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[288\]
+ sky130_fd_sc_hd__dfrtp_1
X_11796_ clknet_leaf_30_clk _00007_ net1201 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07276__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10747_ clknet_leaf_25_clk _00259_ net1185 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[219\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10280__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09017__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10678_ clknet_leaf_59_clk _00190_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[150\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09779__C_N net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06236__C1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06787__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06025__A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09725__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ net808 _02943_ _02944_ net794 vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_121_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10954__RESET_B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10099__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ core.pc.current_pc\[25\] _04591_ net596 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08894__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05722_ _01825_ _01826_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09490_ _05010_ net324 net264 net1774 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a22o_1
XANTENNA__05803__S net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _04528_ _04522_ net228 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05653_ core.register_file.registers_state\[534\] net707 net645 _01757_ vssd1 vssd1
+ vccd1 vccd1 _01758_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08372_ _04451_ _04455_ _04464_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o211a_1
X_05584_ core.register_file.registers_state\[283\] core.register_file.registers_state\[315\]
+ core.register_file.registers_state\[411\] core.register_file.registers_state\[443\]
+ net696 net1012 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_22_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload76_A clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07323_ core.register_file.registers_state\[27\] core.register_file.registers_state\[59\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10271__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07254_ net828 _03357_ _03358_ net977 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08415__A _01958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09008__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06205_ net1045 core.register_file.registers_state\[742\] net750 _02309_ net924 vssd1
+ vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_76_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10985__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07185_ _03289_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout304_A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1046_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06136_ net555 net536 _02208_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06067_ net1025 _02170_ _02171_ net932 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1213_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
Xfanout412 net415 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09716__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 net426 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_8
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
XANTENNA__07727__C1 _03829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout673_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 net458 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_4
Xfanout467 _04667_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_4
X_09826_ _04890_ net2491 net379 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
Xfanout478 net481 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout489 _02487_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_4
XANTENNA__09680__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05753__A1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _04983_ net286 net257 net1633 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06969_ core.register_file.registers_state\[298\] core.register_file.registers_state\[266\]
+ core.register_file.registers_state\[426\] core.register_file.registers_state\[394\]
+ net834 net1069 vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux4_1
XANTENNA__11610__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ net727 _04064_ net525 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ _04887_ net2312 net278 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__mux2_1
XANTENNA__09495__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05505__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07050__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ net462 _04711_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__nand2_2
XANTENNA__05398__D_N net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__B1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11650_ clknet_leaf_49_clk _01162_ net1309 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ clknet_leaf_38_clk _00113_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07258__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11581_ clknet_leaf_31_clk _01093_ net1200 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10262__B1 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10532_ clknet_leaf_76_clk _00044_ net1261 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08207__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10463_ net1380 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10014__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11412__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input67_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10394_ net1392 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07430__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09707__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05441__B1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05684__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10708__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ clknet_leaf_93_clk _00527_ net1239 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08995__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 net993 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08059__X _04164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09486__A2 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07404__A _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07497__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08694__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07497__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08219__B _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07898__X _04003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11848_ clknet_leaf_28_clk net43 net1194 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09238__A2 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11779_ clknet_leaf_24_clk _01283_ net1183 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload11 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_114_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload22 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload22/X sky130_fd_sc_hd__clkbuf_8
Xclkload33 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__inv_6
Xclkload44 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_6
XANTENNA__09946__A0 core.IO_mod.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload55 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_109_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload66 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_8
XFILLER_0_51_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload77 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_8
Xclkload88 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_71_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload99 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_71_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07421__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06855__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07421__B2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ net2512 net429 _04966_ net1000 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05432__B1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ _03083_ _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11633__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07872_ net1113 _03975_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09713__A3 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10005__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09611_ _04978_ net398 net391 net2154 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06823_ _02926_ _02927_ net789 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_69_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06754_ _02857_ _02858_ net792 vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__o21ai_1
X_09542_ _04887_ net2438 net306 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__mux2_1
XANTENNA__09477__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08134__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05705_ net962 _01808_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__or3_1
XANTENNA__07488__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06685_ net1093 core.register_file.registers_state\[851\] core.register_file.registers_state\[883\]
+ net833 net978 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09473_ _04977_ net319 net262 net1923 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_90_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08424_ _01927_ _04491_ _04506_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06696__C1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05636_ net1040 core.register_file.registers_state\[343\] core.register_file.registers_state\[375\]
+ net671 net922 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__o221a_1
XANTENNA__08844__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09229__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08355_ core.pc.current_pc\[12\] _03023_ net576 vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__mux2_1
X_05567_ net638 _01668_ _01669_ _01670_ _01671_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1163_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ _02848_ _02906_ _03409_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07335__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload5 clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_6
XANTENNA__05769__A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06448__C1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08286_ _02277_ _04385_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__nor2_1
X_05498_ net966 _01601_ _01602_ net1006 _01600_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__o311a_1
XFILLER_0_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07237_ net974 _03338_ _03341_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06463__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11163__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__A0 core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ net995 core.register_file.registers_state\[451\] net885 core.register_file.registers_state\[483\]
+ net983 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout790_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout888_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06119_ net1046 core.register_file.registers_state\[584\] core.register_file.registers_state\[616\]
+ net677 net641 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__o221a_1
X_07099_ _03200_ _03203_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1216_X net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07963__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06620__C1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1207 net1208 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10876__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1218 net1224 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_2
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
XANTENNA__05974__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 _04333_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1229 net1236 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_2
XANTENNA__05974__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 _04880_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
Xfanout253 _04683_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout264 _05059_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05791__X _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout275 _05083_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07715__A2 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout286 net288 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_4
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
X_09809_ _05042_ net458 net270 net1886 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06923__B1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08039__B _04016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06687__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11702_ clknet_leaf_71_clk net1588 net1274 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11633_ clknet_leaf_71_clk _01145_ net1274 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05679__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ clknet_leaf_26_clk _01076_ net1203 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ clknet_leaf_36_clk _00027_ net1222 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10250__A3 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11495_ clknet_leaf_65_clk _01007_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[967\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09928__A0 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__A _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10446_ net1416 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10377_ net1430 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06611__C1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10680__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09614__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__B2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08116__C1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09459__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06390__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11036__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
X_06470_ net1034 core.register_file.registers_state\[856\] core.register_file.registers_state\[888\]
+ net666 net923 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08891__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05421_ net655 _01520_ net617 _01519_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__o211ai_1
XANTENNA__08419__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08140_ _04017_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__or2_1
XANTENNA__11186__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05352_ _01388_ _01390_ _01393_ _01395_ net1096 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__o221a_4
XANTENNA__09092__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09631__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08071_ _02345_ _03231_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__nand2_1
Xclkload100 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__clkinv_8
X_05283_ _01387_ _01389_ _01392_ _01394_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__a22o_1
XANTENNA__09919__A0 core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07022_ core.register_file.registers_state\[520\] core.register_file.registers_state\[552\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05653__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08198__A2 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload39_A clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07309__A _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06602__C1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ net2213 net368 _04955_ net434 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__a22o_1
XANTENNA__06213__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold17 core.register_file.registers_state\[957\] vssd1 vssd1 vccd1 vccd1 net1336
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _02902_ _03410_ _02906_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__a21o_1
Xhold28 core.register_file.registers_state\[966\] vssd1 vssd1 vccd1 vccd1 net1347
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 core.register_file.registers_state\[950\] vssd1 vssd1 vccd1 vccd1 net1358
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _03664_ _03800_ _03807_ _02518_ net514 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout371_A _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout469_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ _02907_ _02908_ _02909_ _02910_ net802 net970 vssd1 vssd1 vccd1 vccd1 _02911_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07786_ _03889_ _03890_ net510 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__mux2_1
XANTENNA__06381__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__C1 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _04846_ net395 net307 net1709 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a22o_1
X_06737_ net538 _01957_ _02811_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11562__Q core.decoder.inst\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout636_A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06669__C1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11529__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ net1109 core.register_file.registers_state\[340\] core.register_file.registers_state\[372\]
+ net859 net984 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__o221a_1
X_09456_ _04946_ net316 net311 net2071 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ core.pc.current_pc\[15\] core.pc.current_pc\[16\] _04477_ vssd1 vssd1 vccd1
+ vccd1 _04498_ sky130_fd_sc_hd__and3_1
X_05619_ net1039 core.register_file.registers_state\[983\] core.register_file.registers_state\[1015\]
+ net670 net1010 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09387_ net2021 net329 net322 _04827_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06599_ net777 _02702_ _02703_ net773 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout1166_X net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08338_ _04408_ _04412_ _04421_ _04423_ _04433_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__o311a_1
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09083__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11004__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ _04370_ _04371_ net598 vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o21a_1
XANTENNA__10232__A3 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__B2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ net23 net902 net796 net2318 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__o22a_1
XANTENNA__06841__C1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ clknet_leaf_105_clk _00792_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[752\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08603__A _04139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10231_ net76 net920 vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__and2_1
XANTENNA__10344__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10162_ net1386 net918 net908 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__a21o_1
XANTENNA__07219__A _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_4
Xfanout1015 net1016 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__buf_4
Xfanout1026 net1033 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_4
X_10093_ _04278_ net591 vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__nand2_1
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
Xfanout1048 net1050 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1059 net1061 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10995_ clknet_leaf_12_clk _00507_ net1172 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[467\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_54_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09310__A1 core.register_file.registers_state\[369\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06124__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06124__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09861__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05883__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ clknet_leaf_31_clk _01128_ net1205 vssd1 vssd1 vccd1 vccd1 core.d_hit sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09074__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07085__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11547_ clknet_leaf_23_clk _01059_ net1184 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1019\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08821__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold509 core.register_file.registers_state\[534\] vssd1 vssd1 vccd1 vccd1 net1828
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08513__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11478_ clknet_leaf_61_clk _00990_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[950\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10429_ net1445 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08232__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07388__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07129__A _03231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06033__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05970_ net958 _02073_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__and3_1
Xhold1209 core.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07640_ net452 _02994_ net444 net501 vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a31o_1
X_07571_ _03674_ _03675_ net498 vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
X_06522_ net1096 core.register_file.registers_state\[605\] core.register_file.registers_state\[637\]
+ net837 net803 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__o221a_1
X_09310_ core.register_file.registers_state\[369\] _04666_ _04708_ vssd1 vssd1 vccd1
+ vccd1 _05048_ sky130_fd_sc_hd__o21a_1
XANTENNA__06115__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06115__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09852__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06453_ net965 _02554_ _02557_ net630 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a211o_1
X_09241_ net558 _04840_ _05036_ net339 net2520 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__a32o_1
XFILLER_0_111_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05404_ net896 _01408_ _01410_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__o21a_2
XFILLER_0_8_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ _04952_ net352 net343 net2104 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__a22o_1
X_06384_ net944 core.register_file.registers_state\[833\] net702 core.register_file.registers_state\[865\]
+ net1017 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__a221o_1
XANTENNA__06208__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08123_ _04226_ _04227_ _03695_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05335_ net1315 net1473 net1778 _01443_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
XANTENNA__07615__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06418__A2 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10214__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08812__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout217_A _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05626__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08054_ net491 _04098_ _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__o21ai_4
X_05266_ core.pc.current_pc\[8\] vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07005_ _03100_ _03103_ _03109_ net968 vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__X _05109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A _01379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A2 _04018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09953__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11557__Q core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05929__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _04838_ net601 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__nor2_1
X_07907_ _04008_ _04010_ net485 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__mux2_1
XANTENNA__08879__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net1121 _04714_ net601 vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__or3_4
XANTENNA_fanout753_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07000__C1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ net529 _03918_ _03919_ _03941_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a31oi_1
XANTENNA__06089__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout920_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ net546 _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09508_ _04753_ net400 net309 net1605 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__a22o_1
XANTENNA__11256__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06106__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10780_ clknet_leaf_39_clk _00292_ net1218 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[252\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07502__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ _04912_ net322 net313 net2042 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__a22o_1
XANTENNA__10339__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06118__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11401_ clknet_leaf_38_clk _00913_ net1213 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[873\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08803__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11332_ clknet_leaf_80_clk _00844_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06814__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10891__RESET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06290__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11263_ clknet_leaf_15_clk _00775_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[735\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10214_ net1127 net1395 net912 _05215_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__a31o_1
XANTENNA__08031__A1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11194_ clknet_leaf_8_clk _00706_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[666\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10145_ _03811_ _05190_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__nand2_1
XANTENNA__07891__B _02747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10076_ _04109_ net557 net590 core.pc.current_pc\[10\] net472 vssd1 vssd1 vccd1 vccd1
+ _05145_ sky130_fd_sc_hd__o221a_1
XANTENNA__06345__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06440__S1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11844__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08067__X _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09295__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10978_ clknet_leaf_78_clk _00490_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[450\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07845__A1 _03763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09330__C net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07845__B2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05856__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09598__A1 _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07058__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08270__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 core.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08270__B2 _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06315__X _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold317 core.register_file.registers_state\[447\] vssd1 vssd1 vccd1 vccd1 net1636
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold328 core.register_file.registers_state\[652\] vssd1 vssd1 vccd1 vccd1 net1647
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11224__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold339 core.register_file.registers_state\[875\] vssd1 vssd1 vccd1 vccd1 net1658
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05820__A1_N net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
Xfanout819 net823 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_4
XANTENNA__08897__B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ core.IO_mod.data_from_mem\[27\] core.IO_mod.input_reg\[27\] net251 vssd1
+ vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__mux2_1
XANTENNA__07230__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _04771_ net383 net270 net1654 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__a22o_1
XANTENNA__11374__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 core.register_file.registers_state\[488\] vssd1 vssd1 vccd1 vccd1 net2325
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 core.register_file.registers_state\[629\] vssd1 vssd1 vccd1 vccd1 net2336
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net731 _04278_ net525 _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a211oi_4
XANTENNA__07208__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1028 core.register_file.registers_state\[379\] vssd1 vssd1 vccd1 vccd1 net2347
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05953_ net1036 core.register_file.registers_state\[205\] core.register_file.registers_state\[237\]
+ net666 net651 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__o221a_1
Xhold1039 core.register_file.registers_state\[110\] vssd1 vssd1 vccd1 vccd1 net2358
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05884_ net585 _01988_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__nor2_1
X_08672_ _04670_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07623_ _03726_ _03727_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_85_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05544__C1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07554_ net450 net549 net442 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or3_2
XANTENNA__08628__A3 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06505_ net784 _02608_ _02609_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07836__A1 _03697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07485_ net1100 core.register_file.registers_state\[735\] core.register_file.registers_state\[767\]
+ net844 net822 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_137_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06209__Y _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_A _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1076_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09224_ net563 _04776_ net416 net339 net1556 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06436_ core.register_file.registers_state\[921\] core.register_file.registers_state\[953\]
+ net712 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06367_ net951 core.register_file.registers_state\[578\] net709 core.register_file.registers_state\[610\]
+ net660 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__a221oi_1
X_09155_ _04918_ net351 net343 net1950 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout501_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1243_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05318_ _01393_ _01430_ _01431_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__or3_1
X_08106_ net506 _03715_ _03761_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__o21a_1
XANTENNA__08153__A _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06298_ _02392_ _02395_ _02402_ net718 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__o211ai_4
X_09086_ net2441 net364 net355 _04759_ vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06272__B1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05249_ core.control_logic.instruction\[3\] vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
X_08037_ _03204_ _03205_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05614__A3 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 core.register_file.registers_state\[894\] vssd1 vssd1 vccd1 vccd1 net2159
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold851 core.register_file.registers_state\[239\] vssd1 vssd1 vccd1 vccd1 net2170
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold862 core.register_file.registers_state\[417\] vssd1 vssd1 vccd1 vccd1 net2181
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09683__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap581 _01629_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_1
Xhold873 core.register_file.registers_state\[349\] vssd1 vssd1 vccd1 vccd1 net2192
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 core.register_file.registers_state\[176\] vssd1 vssd1 vccd1 vccd1 net2203
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold895 core.register_file.registers_state\[169\] vssd1 vssd1 vccd1 vccd1 net2214
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A _01372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06024__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06104__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09988_ net1512 net540 net519 _02514_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__a22o_1
XANTENNA__08600__B _03964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10108__C1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ net572 net217 net737 vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__and3_2
XANTENNA__06401__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05783__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__RESET_B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06327__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ clknet_leaf_60_clk _00413_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[373\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06878__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ clknet_leaf_49_clk _01350_ net1311 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05535__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__A1_N net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10832_ clknet_leaf_104_clk _00344_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[304\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06547__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07232__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ clknet_leaf_111_clk _00275_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[235\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05838__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10694_ clknet_leaf_100_clk _00206_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[166\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11247__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05687__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06263__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11315_ clknet_leaf_98_clk _00827_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08998__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08213__D _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ clknet_leaf_89_clk _00758_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[718\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09201__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11177_ clknet_leaf_16_clk _00689_ net1211 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[649\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06566__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ _05178_ _05179_ net556 vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08307__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ _04200_ net592 vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__nand2_1
XANTENNA__06318__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09622__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05829__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07270_ core.register_file.registers_state\[32\] core.register_file.registers_state\[0\]
+ net859 vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06221_ net947 core.register_file.registers_state\[453\] net703 core.register_file.registers_state\[485\]
+ net927 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__RESET_B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05597__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09069__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06152_ _02252_ _02253_ _02255_ net927 net1029 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__o221a_1
XANTENNA__08243__A1 _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09440__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 core.register_file.registers_state\[1012\] vssd1 vssd1 vccd1 vccd1 net1422
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold114 core.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold125 core.ADR_I\[21\] vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
X_06083_ core.register_file.registers_state\[681\] net677 net656 _02187_ vssd1 vssd1
+ vccd1 vccd1 _02188_ sky130_fd_sc_hd__o211a_1
Xhold136 core.CPU_DAT_I\[24\] vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09991__B2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold147 _01213_ vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _01209_ vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09911_ core.control_logic.instruction\[0\] core.CPU_DAT_O\[0\] net893 vssd1 vssd1
+ vccd1 vccd1 _01064_ sky130_fd_sc_hd__mux2_1
Xhold169 core.CPU_DAT_I\[23\] vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10764__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout605 _04670_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_8
Xfanout616 net617 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_8
X_09842_ net203 net2363 net382 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_4
Xfanout638 net642 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_4
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_2
X_09773_ net603 net204 net287 net257 net1984 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_87_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ net1102 core.register_file.registers_state\[201\] core.register_file.registers_state\[233\]
+ net843 net821 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_87_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout284_A _05081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08724_ net605 _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05936_ net945 core.register_file.registers_state\[78\] net704 core.register_file.registers_state\[110\]
+ net657 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a221o_1
XANTENNA__08847__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ core.IO_mod.input_reg\[3\] net254 net729 vssd1 vssd1 vccd1 vccd1 _04727_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout451_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05867_ net1062 core.register_file.registers_state\[721\] core.register_file.registers_state\[753\]
+ net687 net660 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1193_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07606_ _03709_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08586_ net611 net746 _04652_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__or3b_4
X_05798_ core.register_file.registers_state\[658\] core.register_file.registers_state\[690\]
+ net712 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07537_ net449 net551 net441 net502 vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__o31a_1
XFILLER_0_119_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11570__Q core.decoder.inst\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06891__A _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ net617 _03571_ _03572_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09207_ net604 net203 net353 net423 net1706 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__a32o_1
XFILLER_0_134_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06419_ _02346_ _02521_ _02523_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nand3_2
XANTENNA__07690__C1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07399_ _03500_ _03501_ _03503_ _03502_ net793 net828 vssd1 vssd1 vccd1 vccd1 _03504_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1246_X net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08234__A1 _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ _04894_ net1969 net347 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09069_ net613 _04875_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__and2_1
XANTENNA__06340__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11100_ clknet_leaf_62_clk _00612_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[572\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold670 core.ru.prev_busy vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08611__A _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 core.register_file.registers_state\[493\] vssd1 vssd1 vccd1 vccd1 net2000
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 core.register_file.registers_state\[40\] vssd1 vssd1 vccd1 vccd1 net2011
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A1 _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11031_ clknet_leaf_22_clk _00543_ net1181 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10352__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05970__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11200__RESET_B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11864_ clknet_leaf_52_clk _01333_ net1303 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
XANTENNA__05523__A2 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08058__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06720__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06720__B2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10815_ clknet_leaf_15_clk _00327_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11795_ clknet_leaf_29_clk _01299_ net1196 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06159__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10746_ clknet_leaf_7_clk _00258_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[218\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09670__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10280__A1 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10677_ clknet_leaf_62_clk _00189_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[149\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09599__D_N net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08225__B2 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_clk_X clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__A2 _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__B2 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06787__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11359__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ clknet_leaf_16_clk _00741_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[701\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06770_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nor2_1
XANTENNA__09489__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06976__A _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10099__A1 _04317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08894__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05721_ net582 _01782_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08440_ _04526_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08700__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05652_ net949 core.register_file.registers_state\[566\] net763 vssd1 vssd1 vccd1
+ vccd1 _01757_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08371_ _02053_ _04463_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__nand2_1
X_05583_ net1026 _01676_ _01687_ net722 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__o211a_2
XFILLER_0_4_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07322_ core.register_file.registers_state\[155\] core.register_file.registers_state\[187\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09661__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07253_ net1110 core.register_file.registers_state\[672\] core.register_file.registers_state\[640\]
+ net860 net813 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06570__S0 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06204_ net941 core.register_file.registers_state\[710\] vssd1 vssd1 vccd1 vccd1
+ _02309_ sky130_fd_sc_hd__and2_1
XANTENNA__05683__D1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07184_ _03275_ _03276_ _03288_ net769 vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_76_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10009__Y _05105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06135_ net722 _02227_ _02232_ _02239_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07424__C1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06778__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06778__B2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06066_ net936 core.register_file.registers_state\[842\] net693 core.register_file.registers_state\[874\]
+ net1008 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05986__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05450__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_4
XANTENNA__05450__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 net415 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_4
Xfanout424 net426 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_4
XANTENNA__07727__B1 _03827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net440 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09961__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_2
X_09825_ net206 net2062 net382 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XANTENNA__09192__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout468 _04667_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_6
XANTENNA__05738__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net481 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_4
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _04981_ net286 net257 net1634 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__a22o_1
X_06968_ net802 _03069_ _03068_ net789 vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a211o_1
X_08707_ net1723 net466 net431 _04771_ vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__a22o_1
X_05919_ net951 net765 core.register_file.registers_state\[782\] vssd1 vssd1 vccd1
+ vccd1 _02024_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09687_ _04886_ net2384 net280 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06899_ _03000_ _03001_ _03003_ _03002_ net820 net790 vssd1 vssd1 vccd1 vccd1 _03004_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08638_ _04710_ net559 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__nor2_1
XANTENNA__07050__S1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06163__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08569_ _04633_ _04637_ _04643_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ clknet_leaf_14_clk _00112_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ clknet_leaf_27_clk _01092_ net1197 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08606__A _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09652__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06466__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ clknet_leaf_67_clk _00043_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10347__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08207__A1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10462_ net1390 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__A1 core.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10014__B2 _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10393_ net2452 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09183__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ clknet_leaf_98_clk _00526_ net1160 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[486\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11435__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08995__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_8
Xfanout991 net993 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05904__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07391__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input15_X net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08143__B1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09891__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__B2 _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ clknet_leaf_24_clk net42 net1183 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08446__A1 _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ clknet_leaf_28_clk _01282_ net1196 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09643__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09111__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06457__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ clknet_leaf_38_clk _00241_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[201\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload12 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_114_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload23 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_8
Xclkload34 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_4
Xclkload45 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__09946__A1 core.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05680__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload56 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload67 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_8
Xclkload78 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_110_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload89 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_45_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_53_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08251__A _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06855__S1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05968__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07940_ _03086_ _03115_ _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__or3_1
XANTENNA__11193__RESET_B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09174__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ net1006 net900 net546 _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06607__S1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10005__B _02083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09610_ _04976_ net400 net393 net2102 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__a22o_1
XANTENNA__07724__A3 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06822_ net1092 core.register_file.registers_state\[205\] core.register_file.registers_state\[237\]
+ net831 net816 vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_111_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _04886_ net2357 net304 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__mux2_1
X_06753_ net1111 core.register_file.registers_state\[209\] core.register_file.registers_state\[241\]
+ net857 net827 vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_65_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05704_ net1058 core.register_file.registers_state\[469\] core.register_file.registers_state\[501\]
+ net683 net1019 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__o221a_1
X_09472_ _04975_ net321 net263 net1741 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__a22o_1
XANTENNA__10021__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06684_ net1093 core.register_file.registers_state\[979\] core.register_file.registers_state\[1011\]
+ net833 net1072 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__o221a_1
XANTENNA__09882__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08423_ _01897_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05635_ net959 _01739_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ core.pc.current_pc\[11\] _04449_ net597 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09634__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05566_ net937 core.register_file.registers_state\[699\] net748 net1012 vssd1 vssd1
+ vccd1 vccd1 _01671_ sky130_fd_sc_hd__o211a_1
XANTENNA__05402__X _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10244__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07305_ _03403_ _03407_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08285_ _02277_ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05497_ net1058 core.register_file.registers_state\[860\] core.register_file.registers_state\[892\]
+ net683 net927 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__o221a_1
Xclkload6 clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_8
XFILLER_0_117_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1156_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07236_ net1087 _03339_ _03340_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05671__A1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07167_ net994 core.register_file.registers_state\[323\] net885 core.register_file.registers_state\[355\]
+ net1078 vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06118_ net1046 core.register_file.registers_state\[712\] vssd1 vssd1 vccd1 vccd1
+ _02223_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07098_ _02316_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout783_A _01462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05423__B2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06049_ net616 _02150_ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_54_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__clkbuf_2
Xfanout210 _04865_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1111_X net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1219 net1224 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__clkbuf_4
Xfanout232 _05248_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09691__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1209_X net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09165__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout243 _04875_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
XANTENNA_fanout950_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 _03687_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_4
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_4
X_09808_ _04867_ net390 net272 net1628 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__a22o_1
XANTENNA__10180__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _05080_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
XANTENNA__06384__C1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06923__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__A _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _04950_ net287 net274 net2233 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__a22o_1
XANTENNA__08125__A0 _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ clknet_leaf_76_clk net1466 net1260 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11632_ clknet_leaf_76_clk _01144_ net1260 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05312__X _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08979__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ clknet_leaf_26_clk _01075_ net1191 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10514_ clknet_leaf_37_clk _00026_ net1222 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11494_ clknet_leaf_105_clk _01006_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[966\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_126_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07894__B _02747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ net1342 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05695__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08071__A _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ net1399 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__05414__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05414__B2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10106__A _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10825__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09156__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07167__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10171__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__B2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10975__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06127__C1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09864__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05420_ _01517_ _01518_ net622 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09616__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05351_ net1085 _01397_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09092__B2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08070_ net530 _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__nand2_1
X_05282_ _01388_ _01390_ _01393_ _01395_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__o22a_4
XFILLER_0_125_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07642__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload101 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09919__A1 core.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07021_ net772 _03120_ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__or3_1
XFILLER_0_125_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09077__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09395__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05405__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08972_ net570 net210 net739 vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_90_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09364__X _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ net530 _04007_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09147__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 core.register_file.registers_state\[936\] vssd1 vssd1 vccd1 vccd1 net1337
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 core.register_file.registers_state\[1014\] vssd1 vssd1 vccd1 vccd1 net1348
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07854_ _03908_ _03911_ net494 vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10162__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05708__A2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ core.register_file.registers_state\[525\] core.register_file.registers_state\[557\]
+ net863 vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07785_ _02519_ _03763_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__or2_2
XANTENNA__06381__A2 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09524_ _04711_ _04840_ net456 net307 net1960 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__a32o_1
X_06736_ _02840_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__inv_2
XANTENNA__07044__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09455_ _04944_ net316 net311 net2244 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout531_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06667_ core.register_file.registers_state\[276\] core.register_file.registers_state\[308\]
+ core.register_file.registers_state\[404\] core.register_file.registers_state\[436\]
+ net889 net1080 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__mux4_1
XANTENNA__07330__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07330__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_A _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1273_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ _04494_ _04495_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09870__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05618_ net1039 core.register_file.registers_state\[855\] core.register_file.registers_state\[887\]
+ net670 net922 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__o221a_1
XANTENNA__06375__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09386_ net1913 net329 net324 _04821_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__a22o_1
XANTENNA__07881__A2 _03412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06598_ net783 _02694_ _02697_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08337_ _04408_ _04412_ _04421_ _04423_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_43_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05549_ net922 _01650_ _01651_ _01653_ net958 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout1061_X net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09686__S net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07094__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ core.pc.current_pc\[4\] _04361_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout998_A _01368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05644__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07219_ _03319_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__nand2_1
XANTENNA__06841__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05644__B2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08199_ _03759_ _03773_ _03980_ _03771_ _04303_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08603__B _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10230_ net1127 net1625 net913 _05223_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09386__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06404__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10161_ wb.curr_state\[1\] net1125 wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _05205_
+ sky130_fd_sc_hd__and3b_4
XANTENNA__05947__A2 _02051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1005 net1007 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_6
Xfanout1016 core.decoder.inst\[22\] vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_4
Xfanout1027 net1028 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_4
X_10092_ core.pc.current_pc\[16\] net591 vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1038 net1053 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10360__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05962__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06357__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06372__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08649__A1 core.IO_mod.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05580__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ clknet_leaf_70_clk _00506_ net1275 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09310__A2 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11885__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11615_ clknet_leaf_29_clk _01127_ net1198 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05883__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11623__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09074__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06507__S0 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07085__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11546_ clknet_leaf_6_clk _01058_ net1145 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1018\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07180__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11477_ clknet_leaf_63_clk _00989_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[949\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09377__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ net1321 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07388__A1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10359_ _05111_ net1571 net234 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05494__S0 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06994__S0 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ net451 _03536_ net443 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__and3_2
XFILLER_0_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09837__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06521_ net1096 core.register_file.registers_state\[733\] core.register_file.registers_state\[765\]
+ net837 net823 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09301__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09240_ core.register_file.registers_state\[311\] net474 net544 vssd1 vssd1 vccd1
+ vccd1 _05036_ sky130_fd_sc_hd__o21a_1
XANTENNA__05323__B1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06452_ _02555_ _02556_ net1032 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06520__C1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05403_ core.decoder.inst\[30\] net898 net593 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11555__RESET_B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09171_ _04950_ net352 net343 net1631 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__a22o_1
X_06383_ core.decoder.inst\[8\] _01409_ _01411_ net1028 vssd1 vssd1 vccd1 vccd1 _02488_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_8_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08122_ net514 _04119_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__nand2_1
X_05334_ _01428_ _01440_ _01446_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload51_A clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08053_ net496 _04105_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__or2_1
XANTENNA__06823__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05265_ core.pc.current_pc\[2\] vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08423__B _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07004_ net972 _03107_ _03108_ _03106_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_92_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09368__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07379__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11838__Q core.IO_mod.input_reg\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07379__B2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1021_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06587__C1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08955_ net2316 net369 _04943_ net437 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout579_A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _04010_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__inv_2
XANTENNA__10033__X _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1227_A core.register_file.registers_state\[369\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08886_ core.decoder.inst\[8\] net741 vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_32_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07000__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ net484 _03718_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__nor2_1
XANTENNA__06354__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _01664_ _03476_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _04748_ net397 net308 net1671 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06719_ net1108 core.register_file.registers_state\[466\] core.register_file.registers_state\[498\]
+ net858 net1080 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout913_A _01449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ _02519_ _03789_ _03803_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06106__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09438_ _04910_ net318 net311 net2190 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05865__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05865__B2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ net2295 net330 net323 _04731_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ clknet_leaf_13_clk _00912_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[872\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08173__X _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11225__RESET_B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__A _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05617__A1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10071__C1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11331_ clknet_leaf_66_clk _00843_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09359__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06290__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11262_ clknet_leaf_95_clk _00774_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[734\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11748__Q net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11026__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10213_ net98 net915 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__and2_1
X_11193_ clknet_leaf_68_clk _00705_ net1267 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[665\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07517__X _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _03811_ _05190_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or2_1
XANTENNA__08319__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07790__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10075_ net472 _05143_ _05144_ net517 net1448 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a32o_1
XANTENNA__09531__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06750__C1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09295__A1 _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ clknet_leaf_86_clk _00489_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06309__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09047__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09598__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07153__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11529_ clknet_leaf_38_clk _01041_ net1213 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1001\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_29_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 core.register_file.registers_state\[540\] vssd1 vssd1 vccd1 vccd1 net1626
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06281__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold318 core.register_file.registers_state\[282\] vssd1 vssd1 vccd1 vccd1 net1637
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06281__B2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold329 core.CPU_DAT_I\[15\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10365__A0 _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06979__A _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout809 net811 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07230__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08897__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ core.IO_mod.data_from_mem\[16\] net246 _04798_ vssd1 vssd1 vccd1 vccd1 _04799_
+ sky130_fd_sc_hd__a21oi_4
Xhold1007 core.register_file.registers_state\[373\] vssd1 vssd1 vccd1 vccd1 net2326
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 core.register_file.registers_state\[706\] vssd1 vssd1 vccd1 vccd1 net2337
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05952_ net1036 core.register_file.registers_state\[77\] core.register_file.registers_state\[109\]
+ net665 net636 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__o221a_1
Xhold1029 core.register_file.registers_state\[331\] vssd1 vssd1 vccd1 vccd1 net2348
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10530__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07208__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08671_ net728 _04186_ _04718_ _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a211o_2
XANTENNA__11669__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05883_ net1106 net897 _01867_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07622_ net454 _03231_ net446 net500 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05544__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07553_ _02384_ _03656_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__or2_4
XFILLER_0_53_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06504_ net1101 core.register_file.registers_state\[221\] core.register_file.registers_state\[253\]
+ net845 net821 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07484_ net806 _03587_ _03588_ net1085 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05847__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ _04771_ net416 net339 net1754 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05847__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06435_ _02536_ _02537_ _02538_ _02539_ net624 net648 vssd1 vssd1 vccd1 vccd1 _02540_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09038__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout327_A _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07049__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ _04916_ net355 net344 net1843 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__a22o_1
XANTENNA__09589__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06366_ net634 _02470_ _01511_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11049__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08105_ net500 _03725_ _03766_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__o21ba_1
X_05317_ core.decoder.inst\[12\] core.decoder.inst\[14\] net1005 net1012 vssd1 vssd1
+ vccd1 vccd1 _01431_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09085_ net2243 net365 net358 _04752_ vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__a22o_1
XANTENNA__08261__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06297_ net965 _02396_ _02401_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1236_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06272__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ _03175_ _03176_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold830 core.register_file.registers_state\[587\] vssd1 vssd1 vccd1 vccd1 net2149
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10689__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold841 core.register_file.registers_state\[478\] vssd1 vssd1 vccd1 vccd1 net2160
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 core.register_file.registers_state\[847\] vssd1 vssd1 vccd1 vccd1 net2171
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold863 core.register_file.registers_state\[61\] vssd1 vssd1 vccd1 vccd1 net2182
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold874 core.register_file.registers_state\[887\] vssd1 vssd1 vccd1 vccd1 net2193
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1024_X net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 core.register_file.registers_state\[243\] vssd1 vssd1 vccd1 vccd1 net2204
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 core.register_file.registers_state\[468\] vssd1 vssd1 vccd1 vccd1 net2215
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06024__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09761__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ net1804 net542 net521 _02451_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__A1 core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__C _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08938_ net217 net737 vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__and2_1
XANTENNA__10108__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _04655_ _04826_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nor2_2
XFILLER_0_93_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ clknet_leaf_51_clk _00412_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[372\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11880_ clknet_leaf_70_clk _01349_ net1276 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06732__C1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__A _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07513__A _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ clknet_leaf_83_clk _00343_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[303\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09277__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10762_ clknet_leaf_111_clk _00274_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[234\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05838__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09029__B2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ clknet_leaf_96_clk _00205_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[165\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07659__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06416__X _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06135__Y _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11314_ clknet_leaf_67_clk _00826_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10347__A0 _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11245_ clknet_leaf_3_clk _00757_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[717\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09201__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09752__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11176_ clknet_leaf_12_clk _00688_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09606__C net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10127_ core.pc.current_pc\[27\] _05172_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05774__B1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06971__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10058_ core.pc.current_pc\[3\] net591 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__or2_1
XANTENNA__06318__A2 _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09114__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09268__A1 _04887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11147__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08806__X _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06220_ net947 core.register_file.registers_state\[325\] net703 core.register_file.registers_state\[357\]
+ net1017 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06151_ core.register_file.registers_state\[295\] core.register_file.registers_state\[263\]
+ core.register_file.registers_state\[423\] core.register_file.registers_state\[391\]
+ net682 net1017 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09069__B _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold104 core.register_file.registers_state\[20\] vssd1 vssd1 vccd1 vccd1 net1423
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 core.register_file.registers_state\[962\] vssd1 vssd1 vccd1 vccd1 net1434
+ sky130_fd_sc_hd__dlygate4sd3_1
X_06082_ net1051 core.register_file.registers_state\[649\] vssd1 vssd1 vccd1 vccd1
+ _02187_ sky130_fd_sc_hd__or2_1
Xhold126 core.register_file.registers_state\[955\] vssd1 vssd1 vccd1 vccd1 net1445
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _01225_ vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 net153 vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold159 core.ADR_I\[27\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09910_ net1116 _05021_ net461 net377 net1914 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_74_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10338__A0 _02451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06006__A1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout606 _04669_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_4
X_09841_ _04865_ net2391 net381 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
Xfanout617 _01524_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_6
XANTENNA__07203__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09743__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout628 _01522_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_6
Xfanout639 net642 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_4
XANTENNA__11491__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _05012_ net287 net257 net1858 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__a22o_1
X_06984_ net1102 core.register_file.registers_state\[73\] core.register_file.registers_state\[105\]
+ net843 net806 vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_87_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ net727 _04074_ net525 _04784_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a211o_2
X_05935_ _02037_ _02039_ net618 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout277_A _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ net1964 net468 net438 _04726_ vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05866_ _01969_ _01970_ net1031 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__o21a_1
XANTENNA__06714__C1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07605_ net453 _02931_ net445 net502 vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11570__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ _04654_ net615 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__nand2_2
XFILLER_0_135_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05797_ core.register_file.registers_state\[530\] net692 net662 _01901_ vssd1 vssd1
+ vccd1 vccd1 _01902_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1186_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07536_ net449 net551 net441 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__or3_1
XANTENNA__09959__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07809__A2 _03909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08863__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07467_ net1055 core.register_file.registers_state\[223\] core.register_file.registers_state\[255\]
+ net683 net659 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09206_ _05015_ net355 net424 net1799 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__a22o_1
XANTENNA__06493__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06418_ net554 _02273_ _02275_ _02316_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__o211a_2
XFILLER_0_9_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07398_ core.register_file.registers_state\[921\] core.register_file.registers_state\[953\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09137_ _04893_ net1849 net347 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__mux2_1
X_06349_ _01506_ _02451_ _02452_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__o21a_1
XANTENNA__08234__A2 _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06245__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09694__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_X net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09982__A2 _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ net2388 net427 _05017_ net435 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout980_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05453__C1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06340__S1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ _03397_ _03399_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11834__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold660 core.register_file.registers_state\[35\] vssd1 vssd1 vccd1 vccd1 net1979
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 core.register_file.registers_state\[325\] vssd1 vssd1 vccd1 vccd1 net1990
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08611__B _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11030_ clknet_leaf_58_clk _00542_ net1287 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[502\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold682 core.register_file.registers_state\[86\] vssd1 vssd1 vccd1 vccd1 net2001
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07067__X _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold693 core.register_file.registers_state\[818\] vssd1 vssd1 vccd1 vccd1 net2012
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08170__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ clknet_leaf_50_clk _01332_ net1308 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11214__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06181__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10814_ clknet_leaf_93_clk _00326_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[286\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11240__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11794_ clknet_leaf_29_clk _01298_ net1196 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06159__S1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10745_ clknet_leaf_54_clk _00257_ net1299 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[217\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10280__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10676_ clknet_leaf_55_clk _00188_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[148\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05692__C1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06236__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06025__C net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05995__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09186__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ clknet_leaf_41_clk _00740_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[700\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07197__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ clknet_leaf_22_clk _00671_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06944__C1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire245_A _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__X _03810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10099__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05720_ _01811_ _01823_ net587 _01805_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08697__C1 _04762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08161__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05651_ net659 _01754_ _01755_ net962 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_67_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08370_ _02053_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or2_1
X_05582_ _01681_ _01686_ net959 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07347__S0 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07321_ core.register_file.registers_state\[219\] core.register_file.registers_state\[251\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09661__A1 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10271__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07252_ core.register_file.registers_state\[544\] core.register_file.registers_state\[512\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__mux2_1
XANTENNA__05401__A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06203_ net1045 core.register_file.registers_state\[614\] net750 _02307_ vssd1 vssd1
+ vccd1 vccd1 _02308_ sky130_fd_sc_hd__a31o_1
XANTENNA__06570__S1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09413__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07183_ net781 _03285_ _03287_ net967 vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06134_ net632 _02235_ _02238_ net717 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__o31a_1
XFILLER_0_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08712__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05435__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06065_ net936 core.register_file.registers_state\[970\] net693 core.register_file.registers_state\[1002\]
+ net923 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09716__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout403 net404 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_2
XANTENNA__11846__Q core.IO_mod.input_reg\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07727__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__Y _05113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout425 net426 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_6
XANTENNA_fanout394_A _05066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 net440 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_4
Xfanout447 net448 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_2
X_09824_ net222 net2397 net379 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1101_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 _05060_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08858__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06935__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout469 _04667_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_2
XFILLER_0_119_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06967_ _03070_ _03071_ net784 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _04979_ net290 net257 net1680 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout561_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net563 _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__and2_1
X_05918_ net1062 core.register_file.registers_state\[814\] net754 vssd1 vssd1 vccd1
+ vccd1 _02023_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11069__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ _04885_ net1838 net279 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__mux2_1
X_06898_ core.register_file.registers_state\[588\] core.register_file.registers_state\[620\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08637_ net1117 _04660_ _04661_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11581__Q core.decoder.inst\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05849_ _01952_ _01953_ net1027 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10201__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06163__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_X net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A _01459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07360__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09689__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ _04633_ _04637_ _04643_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09101__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07519_ _03619_ net548 _03623_ _03616_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nor4b_4
XTAP_TAPCELL_ROW_61_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ net1124 net596 _04581_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08606__B _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10530_ clknet_leaf_77_clk _00042_ net1262 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06466__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05311__A core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10461_ net1501 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08207__A2 _01395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06218__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10014__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ net1372 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08622__A _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05426__C1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10363__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05977__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09168__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 core.register_file.registers_state\[359\] vssd1 vssd1 vccd1 vccd1 net1809
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11013_ clknet_leaf_92_clk _00525_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[485\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07525__X _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net973 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_4
Xfanout981 _01370_ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10604__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08143__A1 _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1190 core.register_file.registers_state\[375\] vssd1 vssd1 vccd1 vccd1 net2509
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06154__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10111__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ clknet_leaf_37_clk net41 net1223 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08446__A2 _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11777_ clknet_leaf_29_clk _01281_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09643__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06457__A1 core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ clknet_leaf_14_clk _00240_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[200\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10659_ clknet_leaf_67_clk _00171_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[131\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload13 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__bufinv_16
Xclkload24 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_4
XFILLER_0_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload35 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__inv_6
Xclkload46 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_16
XANTENNA__05680__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload57 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_6
XFILLER_0_80_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07957__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload68 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_110_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload79 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_80_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09159__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05432__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _01746_ net552 vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06821_ net1091 core.register_file.registers_state\[77\] core.register_file.registers_state\[109\]
+ net831 net802 vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_108_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ _04885_ net1880 net303 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06752_ net1111 core.register_file.registers_state\[81\] core.register_file.registers_state\[113\]
+ net857 net812 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05703_ net1056 core.register_file.registers_state\[341\] core.register_file.registers_state\[373\]
+ net684 net928 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__o221a_1
X_09471_ _04973_ net320 net262 net2054 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a22o_1
X_06683_ net1084 _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__or2_1
XANTENNA__09882__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08422_ core.pc.current_pc\[18\] _02841_ net576 vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06696__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05634_ core.register_file.registers_state\[279\] core.register_file.registers_state\[311\]
+ core.register_file.registers_state\[407\] core.register_file.registers_state\[439\]
+ net716 net1011 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06696__B2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload81_A clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _04440_ _04441_ _04448_ net209 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a2bb2o_1
X_05565_ net1041 net748 core.register_file.registers_state\[667\] vssd1 vssd1 vccd1
+ vccd1 _01670_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07304_ _02902_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06448__A1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ core.pc.current_pc\[6\] _03200_ net576 vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05496_ net1058 core.register_file.registers_state\[988\] core.register_file.registers_state\[1020\]
+ net683 net1024 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload7/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__07740__S0 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07235_ net990 core.register_file.registers_state\[449\] net875 core.register_file.registers_state\[481\]
+ net982 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1051_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1149_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ core.register_file.registers_state\[291\] core.register_file.registers_state\[259\]
+ core.register_file.registers_state\[419\] core.register_file.registers_state\[387\]
+ net857 net1078 vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07948__B2 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06117_ net942 core.register_file.registers_state\[744\] net761 vssd1 vssd1 vccd1
+ vccd1 _02222_ sky130_fd_sc_hd__or3_1
X_07097_ net538 _02522_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__nand2_1
XANTENNA__05959__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06620__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06048_ net620 _02151_ _02152_ net631 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a31o_1
XANTENNA__06620__B2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11576__Q core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout776_A _01463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 net1314 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout211 _04849_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout222 _04775_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_2
Xfanout233 _05248_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout255 _03734_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1104_X net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06908__C1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout266 net269 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_6
XANTENNA__09570__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 _05083_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_4
X_09807_ net559 _04862_ net456 net270 net2542 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__a32o_1
Xfanout288 _05080_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
X_07999_ _03688_ _04100_ _04101_ net547 _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__o221a_1
Xfanout299 net302 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06384__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ _04948_ net297 net277 net1980 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09322__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08676__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ _04833_ net296 net284 net1894 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07333__C1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ clknet_leaf_76_clk net1668 net1260 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06687__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06687__B2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05895__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ clknet_leaf_76_clk _01143_ net1260 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10358__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09625__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11562_ clknet_leaf_26_clk _01074_ net1203 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05679__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06137__A _02206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ clknet_leaf_46_clk _00025_ net1289 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11493_ clknet_leaf_86_clk _01005_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[965\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05976__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_clk_X clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09389__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ net1360 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07939__A1 _03397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10375_ net1408 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08071__B _03231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06611__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08364__A1 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09614__C net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08116__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09864__A1 _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09122__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11829_ clknet_leaf_49_clk _01330_ net1310 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09616__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08246__B _04350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05350_ net972 net896 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__nor2_2
XFILLER_0_138_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09092__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05281_ _01393_ _01395_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__nor2_1
Xclkload102 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__inv_6
XFILLER_0_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07020_ net1084 _03121_ _03124_ net780 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__o211a_1
XANTENNA__05886__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05653__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06602__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06602__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ net210 net739 vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__and2_1
XANTENNA__06213__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05810__C1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ _03658_ _03731_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__o21bai_2
Xhold19 core.register_file.registers_state\[995\] vssd1 vssd1 vccd1 vccd1 net1338
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08355__A1 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ net493 net265 _03903_ _03956_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a31o_1
XANTENNA__10303__Y _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06366__B1 _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ core.register_file.registers_state\[653\] core.register_file.registers_state\[685\]
+ net863 vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__mux2_1
X_07784_ _03887_ _03888_ net496 vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__mux2_2
XFILLER_0_127_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09304__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06735_ _02827_ _02839_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__nand2_8
X_09523_ _04834_ net401 net310 net1873 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout357_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _04942_ net325 net313 net2266 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__a22o_1
XANTENNA__06669__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06669__B2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06666_ net828 _02767_ _02766_ net787 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__o211a_1
XANTENNA__06656__S net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08405_ _04470_ _04475_ _04484_ _04494_ _04482_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__o311a_1
X_05617_ net1004 _01718_ _01721_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ net1897 net328 net318 _04816_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06597_ _02698_ _02699_ _02701_ _02700_ net786 net810 vssd1 vssd1 vccd1 vccd1 _02702_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09607__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1266_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__nor2_1
XANTENNA__09967__S net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05548_ net938 core.register_file.registers_state\[762\] net757 _01652_ net1010 vssd1
+ vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__o311a_1
XANTENNA__08871__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09083__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07094__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08267_ core.pc.current_pc\[2\] core.pc.current_pc\[3\] core.pc.current_pc\[4\] vssd1
+ vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__and3_1
X_05479_ core.decoder.inst\[28\] net898 net593 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1054_X net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ net494 _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05796__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06841__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08198_ _03788_ _03797_ _04300_ _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout893_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07149_ core.register_file.registers_state\[804\] core.register_file.registers_state\[772\]
+ net854 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10160_ net100 net910 _01450_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__o21a_1
XANTENNA__08610__C_N _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09791__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08900__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_4
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10091_ net473 _05153_ _05154_ net518 net1424 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__a32o_1
Xfanout1017 net1019 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_4
Xfanout1028 net1033 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_4
XANTENNA__08346__A1 _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A0 _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1039 net1041 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07516__A _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__A1 _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06420__A _02146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06357__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08649__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__A1 _04899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ clknet_leaf_73_clk _00505_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08347__A _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05868__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07609__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11614_ clknet_leaf_27_clk _01126_ net1198 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05883__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09074__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06507__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07085__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08282__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11545_ clknet_leaf_60_clk _01057_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1017\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08821__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_67_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07180__S1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11476_ clknet_leaf_56_clk _00988_ net1294 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[948\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_110_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ net1349 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10117__A _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09782__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ _05110_ net2549 net235 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__mux2_1
XANTENNA__06033__C net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05494__S1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ net11 net904 net797 net2455 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__a22o_1
XANTENNA__09534__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09117__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06994__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05571__A1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06520_ net803 _02623_ _02624_ net1085 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05859__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11448__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06451_ net1064 core.register_file.registers_state\[473\] core.register_file.registers_state\[505\]
+ net690 net1022 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05402_ core.decoder.inst\[31\] _01412_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__and2_2
XFILLER_0_17_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09170_ _04948_ net360 net346 net2292 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06382_ net587 _02485_ _02456_ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08121_ net487 _04183_ _04225_ net514 vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__a211o_1
X_05333_ net1129 core.ru.state\[0\] _01441_ _01445_ net893 vssd1 vssd1 vccd1 vccd1
+ _01446_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08273__B1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08812__A2 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10080__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08052_ net528 _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_96_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05264_ net1 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06505__A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ net1101 core.register_file.registers_state\[713\] core.register_file.registers_state\[745\]
+ net845 net821 vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10027__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09773__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08954_ net570 net213 net739 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__and3_1
XANTENNA__06682__S0 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08328__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1014_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09525__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _03633_ _03637_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__and2b_1
XANTENNA__11854__Q core.IO_mod.input_reg\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08885_ core.decoder.inst\[7\] core.decoder.inst\[8\] _01410_ vssd1 vssd1 vccd1 vccd1
+ _04896_ sky130_fd_sc_hd__and3_1
XANTENNA__06339__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07000__A1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07836_ _03697_ _03923_ _03936_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_32_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08866__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07767_ net492 _03870_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout641_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09506_ _04743_ net399 net308 net1772 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__a22o_1
XANTENNA__07839__B1 _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06718_ net1088 _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__or2_1
X_07698_ net451 _02630_ net443 net505 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_45_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07071__A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06649_ net1109 core.register_file.registers_state\[724\] core.register_file.registers_state\[756\]
+ net859 net828 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__o221a_1
X_09437_ _04908_ net321 net313 net2089 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06511__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout906_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_X net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09697__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ net1802 net330 net323 _04725_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07067__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ core.pc.current_pc\[9\] _04413_ net229 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09299_ _04911_ net417 net331 net2037 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08803__A2 _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08614__B _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10071__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ clknet_leaf_79_clk _00842_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06814__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06814__B2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11261_ clknet_leaf_19_clk _00773_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[733\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10965__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10212_ net1128 net1552 net913 _05214_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__a31o_1
XANTENNA__09764__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ clknet_leaf_3_clk _00704_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06578__B1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ net470 _05189_ _05192_ net515 net1977 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09516__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _04123_ net590 vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__nand2_1
XANTENNA_input35_A gpio_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__Q core.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06750__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10976_ clknet_leaf_51_clk _00488_ net1304 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[448\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09295__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05856__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09047__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09400__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07058__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_104_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07153__S1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05608__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11528_ clknet_leaf_9_clk _01040_ net1153 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1000\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06325__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold308 core.ADR_I\[2\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold319 core.register_file.registers_state\[525\] vssd1 vssd1 vccd1 vccd1 net1638
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11890__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11459_ clknet_leaf_65_clk _00971_ net1245 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[931\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09755__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06612__X _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07230__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11120__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07156__A _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09507__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 core.register_file.registers_state\[464\] vssd1 vssd1 vccd1 vccd1 net2327
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05951_ core.register_file.registers_state\[13\] net668 net652 _02055_ vssd1 vssd1
+ vccd1 vccd1 _02056_ sky130_fd_sc_hd__a211o_1
Xhold1019 core.register_file.registers_state\[707\] vssd1 vssd1 vccd1 vccd1 net2338
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08670_ core.IO_mod.data_from_mem\[5\] net246 _04739_ vssd1 vssd1 vccd1 vccd1 _04740_
+ sky130_fd_sc_hd__a21oi_4
X_05882_ net554 _01978_ _01985_ _01986_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__o31a_2
XANTENNA__06995__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ net454 _03260_ net446 net507 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__a31o_1
XANTENNA__05544__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ _02384_ _03656_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nor2_4
XFILLER_0_18_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08089__A3 _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06503_ net1101 core.register_file.registers_state\[93\] core.register_file.registers_state\[125\]
+ net845 net806 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07297__A1 _03397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07483_ net988 core.register_file.registers_state\[703\] net873 core.register_file.registers_state\[671\]
+ net822 vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06434_ core.register_file.registers_state\[601\] core.register_file.registers_state\[633\]
+ net712 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__mux2_1
X_09222_ _04765_ net417 net340 net1787 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09038__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07049__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09153_ _04914_ net355 net344 net2098 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__a22o_1
X_06365_ _02465_ _02469_ _02468_ net964 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10988__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout222_A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08104_ _03386_ _04204_ _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_20_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05316_ core.decoder.inst\[30\] core.decoder.inst\[31\] core.decoder.inst\[7\] net987
+ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_20_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09084_ net2445 net364 net354 _04747_ vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__a22o_1
XANTENNA__09994__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06296_ net1031 _02398_ _02400_ net630 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08153__C _04215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08035_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold820 core.register_file.registers_state\[637\] vssd1 vssd1 vccd1 vccd1 net2139
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1131_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09746__A0 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 core.register_file.registers_state\[355\] vssd1 vssd1 vccd1 vccd1 net2150
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07765__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1229_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold842 core.register_file.registers_state\[611\] vssd1 vssd1 vccd1 vccd1 net2161
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold853 core.register_file.registers_state\[735\] vssd1 vssd1 vccd1 vccd1 net2172
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold864 core.register_file.registers_state\[878\] vssd1 vssd1 vccd1 vccd1 net2183
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 core.register_file.registers_state\[240\] vssd1 vssd1 vccd1 vccd1 net2194
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout689_A _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold886 core.register_file.registers_state\[49\] vssd1 vssd1 vccd1 vccd1 net2205
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 core.register_file.registers_state\[702\] vssd1 vssd1 vccd1 vccd1 net2216
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ _05096_ core.ru.state\[5\] _01447_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__nor3b_1
XANTENNA__06241__Y _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10108__A1 _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ net2340 net367 _04931_ net431 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__a22o_1
XANTENNA__05783__A1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05783__B2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ _04820_ net2498 net374 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07819_ net493 _03853_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__or2_1
XANTENNA__05535__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08799_ net733 _03944_ net526 _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o211a_4
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06732__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08609__B _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10830_ clknet_leaf_86_clk _00342_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[302\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10761_ clknet_leaf_38_clk _00273_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[233\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09029__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10692_ clknet_leaf_77_clk _00204_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[164\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08625__A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05601__X _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10366__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06145__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11313_ clknet_leaf_81_clk _00825_ net1255 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[785\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11143__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05471__B1 _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ clknet_leaf_101_clk _00756_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[716\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09737__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09201__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07212__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ clknet_leaf_91_clk _00687_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10126_ net1124 core.pc.current_pc\[25\] core.pc.current_pc\[26\] core.pc.current_pc\[27\]
+ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__o211a_1
XANTENNA__11293__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10057_ net473 _05132_ _05133_ net517 net1627 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06318__A3 _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09622__C net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10130__A _03964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10959_ clknet_leaf_83_clk _00471_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[431\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10283__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09130__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11187__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06150_ net1055 core.register_file.registers_state\[487\] net753 _02254_ vssd1 vssd1
+ vccd1 vccd1 _02255_ sky130_fd_sc_hd__a31o_1
XANTENNA__08822__X _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09440__A2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold105 core.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06081_ core.register_file.registers_state\[521\] core.register_file.registers_state\[553\]
+ net701 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_1
Xhold116 core.ADR_I\[26\] vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 core.register_file.registers_state\[11\] vssd1 vssd1 vccd1 vccd1 net1446
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05462__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold138 core.register_file.registers_state\[1015\] vssd1 vssd1 vccd1 vccd1 net1457
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 core.register_file.registers_state\[2\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ net204 net2485 net379 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__mux2_1
Xfanout607 _04669_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
Xfanout618 _01524_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout629 _01522_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09771_ _05010_ net297 net259 net1758 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__a22o_1
X_06983_ core.register_file.registers_state\[9\] core.register_file.registers_state\[41\]
+ core.register_file.registers_state\[137\] core.register_file.registers_state\[169\]
+ net872 net821 vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ core.IO_mod.data_from_mem\[13\] net246 _04783_ vssd1 vssd1 vccd1 vccd1 _04784_
+ sky130_fd_sc_hd__a21oi_1
X_05934_ core.register_file.registers_state\[14\] net704 net643 _02038_ vssd1 vssd1
+ vccd1 vccd1 _02039_ sky130_fd_sc_hd__o211a_1
XANTENNA__07614__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09900__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08653_ net572 net608 net225 vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_1_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05865_ net1061 core.register_file.registers_state\[465\] core.register_file.registers_state\[497\]
+ net688 net1021 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08429__B _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07604_ net453 _03023_ net445 net508 vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06190__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05796_ net1062 core.register_file.registers_state\[562\] net755 vssd1 vssd1 vccd1
+ vccd1 _01901_ sky130_fd_sc_hd__and3_1
X_08584_ _04656_ _04657_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nand2_4
XFILLER_0_89_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11016__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07535_ net450 _02747_ net442 vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__or3_4
XFILLER_0_7_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1081_A core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout437_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1179_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07466_ net1058 core.register_file.registers_state\[95\] core.register_file.registers_state\[127\]
+ net683 net645 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06417_ _02346_ _02521_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__nand2_1
X_09205_ net603 net204 net352 net423 net1641 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06493__A2 _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07690__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ core.register_file.registers_state\[985\] core.register_file.registers_state\[1017\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10026__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06348_ _01506_ _02451_ _02452_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ _04849_ net2492 net350 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__mux2_1
XANTENNA__11579__Q core.decoder.inst\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ net566 net604 net203 vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__and3_1
X_06279_ net586 net535 _02382_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a21o_4
XFILLER_0_114_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1134_X net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09719__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ net527 _04111_ _04112_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__o31a_2
XFILLER_0_124_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold650 core.register_file.registers_state\[219\] vssd1 vssd1 vccd1 vccd1 net1969
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_A _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 core.register_file.registers_state\[761\] vssd1 vssd1 vccd1 vccd1 net1980
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold672 core.register_file.registers_state\[609\] vssd1 vssd1 vccd1 vccd1 net1991
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 core.register_file.registers_state\[494\] vssd1 vssd1 vccd1 vccd1 net2002
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 core.register_file.registers_state\[639\] vssd1 vssd1 vccd1 vccd1 net2013
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1301_X net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ net1875 net1678 net799 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07524__A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11862_ clknet_leaf_28_clk net59 net1195 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06181__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07811__X _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10813_ clknet_leaf_17_clk _00325_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[285\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11793_ clknet_leaf_29_clk _01297_ net1200 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11509__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10744_ clknet_leaf_5_clk _00256_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[216\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09670__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07681__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10675_ clknet_leaf_97_clk _00187_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[147\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09958__A0 core.IO_mod.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08630__B1 _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11227_ clknet_leaf_19_clk _00739_ net1190 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[699\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11158_ clknet_leaf_44_clk _00670_ net1287 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[630\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06944__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ net1433 net515 _05164_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_125_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11089_ clknet_leaf_74_clk _00601_ net1255 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[561\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09489__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07434__A _03536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11039__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08697__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08161__A2 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05650_ net1057 core.register_file.registers_state\[726\] vssd1 vssd1 vccd1 vccd1
+ _01755_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_67_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07721__X _03826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05581_ net638 _01682_ _01683_ _01685_ net1004 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a311o_1
XFILLER_0_4_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05380__C1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ net1096 core.register_file.registers_state\[475\] core.register_file.registers_state\[507\]
+ net837 net1070 vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07347__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09661__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07251_ net997 core.register_file.registers_state\[704\] net888 core.register_file.registers_state\[736\]
+ net813 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10008__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06202_ net940 core.register_file.registers_state\[582\] vssd1 vssd1 vccd1 vccd1
+ _02307_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05683__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06880__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07182_ net1088 _03279_ _03280_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_76_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06133_ _02236_ _02237_ net626 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07424__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08712__B net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05828__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06064_ net958 _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__and2_1
XANTENNA__06632__C1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05986__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05530__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05986__B2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout404 _05061_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
XANTENNA__10035__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout415 _05054_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07727__A2 _03826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout426 _05028_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
X_09823_ _04889_ core.register_file.registers_state\[842\] net379 vssd1 vssd1 vccd1
+ vccd1 _00882_ sky130_fd_sc_hd__mux2_1
Xfanout437 net440 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout459 _05060_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_4
XANTENNA_fanout387_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _04977_ net287 net260 net2048 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06966_ net986 core.register_file.registers_state\[202\] net862 core.register_file.registers_state\[234\]
+ net802 vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07344__A _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ net605 _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05917_ _02020_ _02021_ net1006 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a21o_1
X_09685_ _04884_ net2246 net281 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__mux2_1
XANTENNA__10041__Y _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06897_ core.register_file.registers_state\[716\] core.register_file.registers_state\[748\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1296_A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ net1116 _04660_ _04661_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a21boi_4
X_05848_ net1044 core.register_file.registers_state\[464\] core.register_file.registers_state\[496\]
+ net673 net1013 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__o221a_1
XANTENNA__08874__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06163__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08567_ _04641_ _04642_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout721_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05779_ net616 _01882_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout819_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07518_ _01490_ _03620_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08498_ _04577_ _04579_ _04580_ net208 net596 vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__o221ai_1
XANTENNA__09652__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10556__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08606__C _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07449_ core.register_file.registers_state\[735\] core.register_file.registers_state\[767\]
+ net699 vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05311__B _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__C1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ net1403 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08903__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09119_ _04887_ net2427 net348 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
X_10391_ net1405 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08622__B _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05977__A1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 core.register_file.registers_state\[284\] vssd1 vssd1 vccd1 vccd1 net1799
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 core.register_file.registers_state\[39\] vssd1 vssd1 vccd1 vccd1 net1810
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ clknet_leaf_75_clk _00524_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[484\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06926__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout971 net973 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_4
Xfanout982 net985 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 net997 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11772__Q core.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_84_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
Xhold1180 core.register_file.registers_state\[160\] vssd1 vssd1 vccd1 vccd1 net2499
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08143__A2 _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1191 core.register_file.registers_state\[376\] vssd1 vssd1 vccd1 vccd1 net2510
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06154__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11845_ clknet_leaf_36_clk net40 net1221 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11776_ clknet_leaf_28_clk _01280_ net1194 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08085__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06457__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10727_ clknet_leaf_93_clk _00239_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08851__A0 _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10658_ clknet_leaf_78_clk _00170_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[130\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08813__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload14 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_114_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload25 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_8
Xclkload36 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_84_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload47 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__inv_8
Xclkload58 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_12
XFILLER_0_23_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10589_ clknet_leaf_16_clk _00101_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[61\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload69 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_6
XANTENNA__07957__A2 _04060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06333__A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05968__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07863__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06917__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06820_ net817 _02923_ _02924_ net784 vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06751_ net827 _02854_ _02855_ net787 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_75_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05702_ net1030 _01806_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__or2_1
X_09470_ _04971_ net318 net262 net2025 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a22o_1
X_06682_ core.register_file.registers_state\[787\] core.register_file.registers_state\[819\]
+ core.register_file.registers_state\[915\] core.register_file.registers_state\[947\]
+ net865 net1073 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux4_1
XANTENNA__07342__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08421_ core.pc.current_pc\[17\] net599 _04509_ _04510_ vssd1 vssd1 vccd1 vccd1 _00025_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05633_ _01734_ _01737_ net631 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05353__C1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08352_ _04446_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__xnor2_1
X_05564_ net1041 net748 core.register_file.registers_state\[539\] vssd1 vssd1 vccd1
+ vccd1 _01669_ sky130_fd_sc_hd__a21o_1
XANTENNA__09095__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06508__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09634__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload74_A clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07303_ _02900_ _02901_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08842__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__A3 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ core.pc.current_pc\[5\] net599 _04383_ _04384_ vssd1 vssd1 vccd1 vccd1 _00013_
+ sky130_fd_sc_hd__o22a_1
X_05495_ net1030 _01599_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__or2_1
XANTENNA__06227__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05656__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__S1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07234_ net989 core.register_file.registers_state\[321\] net875 core.register_file.registers_state\[353\]
+ net1076 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07165_ net812 _03266_ _03265_ net793 vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1044_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A2 _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06116_ net1038 core.register_file.registers_state\[968\] core.register_file.registers_state\[1000\]
+ net672 net1011 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__o221a_1
XANTENNA__06605__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__inv_2
XANTENNA__11857__Q core.IO_mod.input_reg\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06047_ net935 core.register_file.registers_state\[202\] net693 core.register_file.registers_state\[234\]
+ net636 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1211_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout212 _04844_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
Xfanout223 _04736_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout671_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_4
XANTENNA__09570__A1 _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ net558 _04857_ net456 net270 net1607 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 _05082_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_8
XANTENNA__06384__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07998_ _02176_ _03081_ _03618_ _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__a211o_1
Xfanout289 net291 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_4
XANTENNA__10180__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _04946_ net287 net274 net1820 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__a22o_1
XANTENNA__11592__Q core.IO_mod.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06949_ _01632_ _02176_ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout936_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09322__A1 _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06136__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ _04827_ net293 net284 net2162 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__a22o_1
XANTENNA__09873__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08619_ _03839_ _04672_ _04693_ _03862_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net1116 _04654_ net611 net457 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__or4b_4
XANTENNA__08617__B _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05895__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11630_ clknet_leaf_54_clk _01142_ net1299 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09086__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09625__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ clknet_leaf_25_clk _01073_ net1186 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08833__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05647__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10512_ clknet_leaf_46_clk _00024_ net1290 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08192__X _04297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ clknet_leaf_81_clk _01004_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[964\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10443_ net1402 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06424__Y _02529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07249__A _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input65_A gpio_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08061__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11767__Q core.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ net1490 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__05695__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07495__S0 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10171__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net791 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
XANTENNA__05583__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06127__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08808__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09864__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09403__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11828_ clknet_leaf_49_clk _01329_ net1310 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10871__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07088__C1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ clknet_leaf_31_clk net1692 net1201 vssd1 vssd1 vccd1 vccd1 core.ru.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05638__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05280_ core.control_logic.instruction\[6\] core.control_logic.instruction\[5\] net1123
+ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__nand3b_4
XANTENNA__06835__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload103 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__11227__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07159__A _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08830__X _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07260__C1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ net2017 net367 _04953_ net432 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__a22o_1
XANTENNA__09645__Y _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07921_ net265 _04016_ _04024_ _03972_ _04023_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a221o_1
XANTENNA__06350__X _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07012__C1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07852_ net492 _03897_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__nand2_1
XANTENNA__06366__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05407__A core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ net1091 core.register_file.registers_state\[589\] core.register_file.registers_state\[621\]
+ net831 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__o22a_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
X_07783_ _03756_ _03767_ net484 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_48_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09522_ _04828_ net399 net310 net1857 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a22o_1
X_06734_ net967 _02835_ _02838_ net770 _02832_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a311o_2
XFILLER_0_56_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08718__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07866__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09453_ _04940_ net326 net313 net2303 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__a22o_1
X_06665_ _02768_ _02769_ net793 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout252_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08404_ _04470_ _04475_ _04484_ _04482_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__o31a_1
X_05616_ _01713_ _01719_ _01720_ _01712_ net933 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_47_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09384_ net2185 net329 net324 _04811_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a22o_1
X_06596_ core.register_file.registers_state\[854\] core.register_file.registers_state\[886\]
+ net880 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XANTENNA__09607__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ _02147_ _04430_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05547_ net1039 core.register_file.registers_state\[730\] vssd1 vssd1 vccd1 vccd1
+ _01652_ sky130_fd_sc_hd__or2_1
XANTENNA__08815__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout517_A _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1259_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05629__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08266_ _04354_ _04359_ _04367_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__nor3_1
X_05478_ net555 _01582_ _01552_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07094__A2 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06525__X _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07217_ net504 net477 _01632_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a21o_1
XANTENNA__10047__X _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ net1112 _01780_ _02718_ _04301_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07148_ _03249_ _03250_ _03252_ _03251_ net792 net812 vssd1 vssd1 vccd1 vccd1 _03253_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11587__Q core.IO_mod.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10207__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06054__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout886_A _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07251__C1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07079_ core.register_file.registers_state\[870\] core.register_file.registers_state\[838\]
+ net839 vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08900__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10090_ _04028_ net591 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__nand2_1
Xfanout1007 core.decoder.inst\[23\] vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_8
XFILLER_0_22_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1029 net1033 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_4
XANTENNA__07003__C1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06357__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06420__B _02206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05317__A core.decoder.inst\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06109__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992_ clknet_leaf_105_clk _00504_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[464\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10894__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10369__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11613_ clknet_leaf_29_clk _01125_ net1198 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10208__A3 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire410 _05057_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_2
X_11544_ clknet_leaf_4_clk _01056_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1016\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_108_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11475_ clknet_leaf_11_clk _00987_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[947\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08034__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10426_ net1365 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09231__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09782__A1 _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07242__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10357_ _05109_ net1566 net234 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10288_ net10 net905 _05244_ net2533 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__a22o_1
XANTENNA__06348__A1 _01506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05556__C1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06757__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05661__S net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06450_ net1064 core.register_file.registers_state\[345\] core.register_file.registers_state\[377\]
+ net690 net930 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06520__A1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10776__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05401_ net898 _01504_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__or2_4
XFILLER_0_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06381_ net586 _02485_ _02456_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05332_ core.ru.state\[4\] core.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__or2_1
X_08120_ _03714_ _03942_ _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06284__B1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05263_ core.WRITE_I vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
X_08051_ _03394_ _04142_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_96_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07481__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07002_ net1101 core.register_file.registers_state\[585\] core.register_file.registers_state\[617\]
+ net845 net807 vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o221a_1
XFILLER_0_109_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_71_clk_X clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__B _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09497__A_N net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09773__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06587__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06587__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07617__A _03201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ net213 net739 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06682__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07904_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08884_ net242 net2423 net373 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07835_ net531 _03939_ _03938_ _03658_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_32_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout467_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07766_ net488 net476 _03790_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_49_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05562__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ _04738_ net400 net309 net1861 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__a22o_1
XANTENNA__07839__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ core.register_file.registers_state\[274\] core.register_file.registers_state\[306\]
+ core.register_file.registers_state\[402\] core.register_file.registers_state\[434\]
+ net889 net1079 vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07697_ _03800_ _03801_ net482 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08167__B _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09436_ _04906_ net323 net314 net2073 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__a22o_1
XANTENNA__08882__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06648_ net1109 core.register_file.registers_state\[596\] core.register_file.registers_state\[628\]
+ net860 net813 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05314__A2 _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08735__X _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06511__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09367_ net2181 net329 net321 _04720_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ net969 _02680_ _02683_ net775 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08318_ core.pc.current_pc\[8\] net597 _04416_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09461__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _04909_ net419 net333 net2022 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10071__A1 _04139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__C _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08249_ core.pc.current_pc\[3\] _03289_ net577 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07472__C1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ clknet_leaf_41_clk _00772_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[732\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08016__B2 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08911__A _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06027__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ net97 net920 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__and2_1
XANTENNA__09764__A1 _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11191_ clknet_leaf_8_clk _00703_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[663\]
+ sky130_fd_sc_hd__dfrtp_1
X_10142_ _05190_ _05191_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__or2_1
XANTENNA__07527__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput190 net190 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_100_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10073_ core.pc.current_pc\[9\] net590 vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or2_1
XANTENNA__11234__RESET_B net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05538__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__Y _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06750__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10975_ clknet_leaf_14_clk _00487_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[447\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05710__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__B net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09452__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06606__A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11527_ clknet_leaf_65_clk _01039_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[999\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold309 core.register_file.registers_state\[828\] vssd1 vssd1 vccd1 vccd1 net1628
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11458_ clknet_leaf_79_clk _00970_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[930\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09204__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10409_ net1350 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__clkbuf_1
X_11389_ clknet_leaf_18_clk _00901_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[861\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06569__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09128__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06341__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05777__C1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05950_ net1037 core.register_file.registers_state\[45\] net747 vssd1 vssd1 vccd1
+ vccd1 _02055_ sky130_fd_sc_hd__and3_1
Xhold1009 core.register_file.registers_state\[163\] vssd1 vssd1 vccd1 vccd1 net2328
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05881_ net586 _01958_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11415__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07620_ net449 _03261_ net441 vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_85_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ _02345_ _03620_ _01492_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__or3b_4
XFILLER_0_92_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06502_ core.register_file.registers_state\[29\] core.register_file.registers_state\[61\]
+ core.register_file.registers_state\[157\] core.register_file.registers_state\[189\]
+ net872 net821 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11565__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09691__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07482_ core.register_file.registers_state\[543\] core.register_file.registers_state\[575\]
+ net873 vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _04760_ net418 net339 net1693 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06433_ core.register_file.registers_state\[537\] core.register_file.registers_state\[569\]
+ net713 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09152_ _04912_ net358 net345 net2250 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__a22o_1
X_06364_ net929 _02467_ net1031 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09443__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08103_ _03618_ _04206_ _04207_ net547 _04205_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__o32a_1
X_05315_ net1114 _01415_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09083_ net2433 net364 net356 _04742_ vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06295_ net1060 core.register_file.registers_state\[483\] net754 _02399_ net929 vssd1
+ vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a311o_1
XANTENNA__09994__B2 _02272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ net528 _04124_ _04136_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_82_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold810 core.register_file.registers_state\[715\] vssd1 vssd1 vccd1 vccd1 net2129
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06009__A0 _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold821 core.register_file.registers_state\[539\] vssd1 vssd1 vccd1 vccd1 net2140
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold832 core.register_file.registers_state\[651\] vssd1 vssd1 vccd1 vccd1 net2151
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07206__C1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold843 core.register_file.registers_state\[693\] vssd1 vssd1 vccd1 vccd1 net2162
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold854 core.register_file.registers_state\[229\] vssd1 vssd1 vccd1 vccd1 net2173
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__B1 _03861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 core.register_file.registers_state\[724\] vssd1 vssd1 vccd1 vccd1 net2184
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 core.register_file.registers_state\[327\] vssd1 vssd1 vccd1 vccd1 net2195
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 core.register_file.registers_state\[443\] vssd1 vssd1 vccd1 vccd1 net2206
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_51_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold898 core.register_file.registers_state\[717\] vssd1 vssd1 vccd1 vccd1 net2217
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ core.ru.state\[0\] net556 _05094_ _05095_ vssd1 vssd1 vccd1 vccd1 _05096_
+ sky130_fd_sc_hd__a211o_4
XANTENNA__06251__A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05768__C1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout584_A _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ net568 net218 net735 vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__and3_1
XANTENNA__08877__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10108__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__X _03739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ net215 net2403 net371 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout751_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__B1 _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07818_ net511 _03922_ _03921_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_19_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08798_ core.IO_mod.data_from_mem\[25\] net247 _04847_ net726 vssd1 vssd1 vccd1 vccd1
+ _04848_ sky130_fd_sc_hd__a211o_1
XANTENNA__06732__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07749_ net489 _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__RESET_B net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09682__A0 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ clknet_leaf_14_clk _00272_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[232\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08906__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10292__A1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09419_ net2215 net214 net408 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XANTENNA__10292__B2 core.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ clknet_leaf_67_clk _00203_ net1268 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[163\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10932__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09434__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11312_ clknet_leaf_104_clk _00824_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[784\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11243_ clknet_leaf_107_clk _00755_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[715\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09201__A3 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__Q core.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ clknet_leaf_99_clk _00686_ net1160 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[646\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _05175_ _05176_ _05092_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__o21ai_1
X_10056_ _04215_ net592 vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07634__A_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08476__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10958_ clknet_leaf_88_clk _00470_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[430\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08476__B2 _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05909__S0 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09411__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10283__B2 core.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10889_ clknet_leaf_38_clk _00401_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[361\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08228__A1 _03739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06080_ net960 _02183_ _02184_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_78_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold106 core.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold117 core.ADR_I\[25\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05998__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05462__A1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold128 core.register_file.registers_state\[25\] vssd1 vssd1 vccd1 vccd1 net1447
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 net182 vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire552_A _02686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__A1 _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout608 net610 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_4
XANTENNA__07203__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11685__Q core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 _01524_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ _05008_ net288 net257 net2317 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__a22o_1
X_06982_ _03056_ _03085_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__and2_1
XANTENNA__10805__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ core.IO_mod.input_reg\[13\] net251 net725 vssd1 vssd1 vccd1 vccd1 _04783_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05933_ net946 core.register_file.registers_state\[46\] net766 vssd1 vssd1 vccd1
+ vccd1 _02038_ sky130_fd_sc_hd__or3_1
Xfanout1190 net1209 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__buf_2
XANTENNA__07614__B _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ net608 net225 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__and2_1
X_05864_ net1060 core.register_file.registers_state\[337\] core.register_file.registers_state\[369\]
+ net688 net929 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_1_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06714__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06714__B2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ _03706_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__nand2_1
X_08583_ _04656_ _04657_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10955__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05922__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05795_ _01898_ _01899_ net1032 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07534_ _03635_ _03638_ net485 vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__mux2_1
XANTENNA__08467__A1 _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09664__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06478__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10274__B2 core.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07465_ _03567_ _03569_ net626 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout332_A _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1074_A core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09204_ _05012_ net353 net423 net1637 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__a22o_1
X_06416_ net504 net492 net477 _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_63_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06246__A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07396_ core.register_file.registers_state\[857\] core.register_file.registers_state\[889\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__mux2_1
XANTENNA__10039__Y _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10026__B2 _05113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09967__A1 core.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07427__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ net212 net2275 net347 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__mux2_1
X_06347_ net554 _02424_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1241_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09066_ net2254 net428 _05016_ net998 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06278_ _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__inv_2
XANTENNA__06245__A3 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05453__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout799_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ _03658_ _03923_ _04116_ _04121_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__o211a_2
XANTENNA__05453__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06650__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 core.register_file.registers_state\[90\] vssd1 vssd1 vccd1 vccd1 net1959
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold651 core.register_file.registers_state\[48\] vssd1 vssd1 vccd1 vccd1 net1970
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold662 core.register_file.registers_state\[508\] vssd1 vssd1 vccd1 vccd1 net1981
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08611__D _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09195__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 core.register_file.registers_state\[422\] vssd1 vssd1 vccd1 vccd1 net1992
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold684 core.register_file.registers_state\[117\] vssd1 vssd1 vccd1 vccd1 net2003
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 core.register_file.registers_state\[360\] vssd1 vssd1 vccd1 vccd1 net2014
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10215__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout966_A _01373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06402__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ net1505 core.CPU_DAT_O\[24\] net798 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__mux2_1
XANTENNA__09292__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ net2229 net367 _04919_ net431 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ net1120 _05076_ net376 net1735 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__a22o_1
XANTENNA__06705__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ clknet_leaf_28_clk net58 net1194 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10812_ clknet_leaf_40_clk _00324_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ clknet_leaf_29_clk _01296_ net1200 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09655__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10743_ clknet_leaf_22_clk _00255_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[215\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10674_ clknet_leaf_71_clk _00186_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08642__Y _04716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07969__B1 _04073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08091__C1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05995__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09186__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ clknet_leaf_9_clk _00738_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[698\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07197__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ clknet_leaf_63_clk _00669_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[629\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06944__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ _03985_ net557 net588 core.pc.current_pc\[23\] net470 vssd1 vssd1 vccd1 vccd1
+ _05164_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_125_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09406__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11088_ clknet_leaf_104_clk _00600_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[560\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10978__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _01502_ _01549_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_121_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09894__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05580_ net937 core.register_file.registers_state\[763\] net748 _01684_ net1010 vssd1
+ vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__o2111a_1
XANTENNA__06765__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05380__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09141__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10256__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07121__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07250_ net996 core.register_file.registers_state\[576\] net888 core.register_file.registers_state\[608\]
+ net828 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07672__A2 _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06201_ net940 core.register_file.registers_state\[646\] net697 core.register_file.registers_state\[678\]
+ net639 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a221o_1
XANTENNA__05683__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10008__B2 _05104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06880__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07181_ net1079 _03278_ _03277_ net976 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11337__RESET_B net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06132_ net1047 core.register_file.registers_state\[200\] core.register_file.registers_state\[232\]
+ net678 net656 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__o221a_1
XFILLER_0_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08281__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05435__B2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06063_ core.register_file.registers_state\[810\] core.register_file.registers_state\[778\]
+ core.register_file.registers_state\[938\] core.register_file.registers_state\[906\]
+ net667 net1008 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05530__S1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout405 net411 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_6
XANTENNA__08385__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout416 net418 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_4
X_09822_ _04888_ net2511 net379 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
Xfanout427 net430 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_8
Xfanout438 net440 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10192__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_2
XANTENNA__07184__X _03289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__RESET_B net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ _04975_ net295 net258 net1650 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__a22o_1
X_06965_ net986 core.register_file.registers_state\[74\] net862 core.register_file.registers_state\[106\]
+ net816 vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ net732 _04767_ _04768_ _04766_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a31o_4
XANTENNA__05416__Y _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05916_ net1054 core.register_file.registers_state\[686\] core.register_file.registers_state\[654\]
+ net681 net644 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a221o_1
XANTENNA__08688__A1 core.IO_mod.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ net223 net1962 net280 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__mux2_1
X_06896_ core.register_file.registers_state\[652\] core.register_file.registers_state\[684\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
XANTENNA__09885__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07912__X _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08635_ net475 net545 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nand2_1
X_05847_ net1044 core.register_file.registers_state\[336\] core.register_file.registers_state\[368\]
+ net673 net924 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout547_A _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07360__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1289_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08566_ _01386_ net549 net574 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05778_ net1046 core.register_file.registers_state\[595\] core.register_file.registers_state\[627\]
+ net676 net637 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__o221a_1
XANTENNA__09637__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07517_ _01500_ _03620_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__or2_4
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09101__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08497_ net1124 _04562_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_X net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07448_ core.register_file.registers_state\[671\] core.register_file.registers_state\[703\]
+ net700 vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06466__A3 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06871__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05311__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11078__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ net1108 core.register_file.registers_state\[473\] core.register_file.registers_state\[505\]
+ net858 net1080 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09118_ _04886_ net2299 net349 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11007__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ net1423 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08622__C _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05426__B2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09049_ net744 net464 _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__and3_1
XANTENNA__07519__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06423__B _01987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09168__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold470 core.register_file.registers_state\[621\] vssd1 vssd1 vccd1 vccd1 net1789
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold481 core.register_file.registers_state\[857\] vssd1 vssd1 vccd1 vccd1 net1800
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 net141 vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ clknet_leaf_73_clk _00523_ net1272 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10183__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net957 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_2
XANTENNA__07535__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout961 _01373_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout972 net973 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08128__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout983 net985 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_4
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1170 core.register_file.registers_state\[142\] vssd1 vssd1 vccd1 vccd1 net2489
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09876__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1181 core.register_file.registers_state\[333\] vssd1 vssd1 vccd1 vccd1 net2500
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09340__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1192 core.register_file.registers_state\[841\] vssd1 vssd1 vccd1 vccd1 net2511
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09891__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ clknet_leaf_29_clk net39 net1195 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09628__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05362__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ clknet_leaf_24_clk _01279_ net1183 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09643__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10726_ clknet_leaf_106_clk _00238_ net1160 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[198\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08653__X _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10657_ clknet_leaf_84_clk _00169_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[129\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08813__B _04860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload15 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_6
Xclkload26 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_4
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload37 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_12
XANTENNA__06614__A _01781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10588_ clknet_leaf_39_clk _00100_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09800__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload48 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload59 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09159__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ clknet_leaf_16_clk _00721_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10174__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06917__A1 _01462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09136__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08119__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06750_ net1111 core.register_file.registers_state\[177\] net856 core.register_file.registers_state\[145\]
+ net812 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09867__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05701_ core.register_file.registers_state\[277\] core.register_file.registers_state\[309\]
+ core.register_file.registers_state\[405\] core.register_file.registers_state\[437\]
+ net707 net1024 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux4_1
X_06681_ _02752_ _02785_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__or2_1
XANTENNA__07342__A1 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ _04502_ _04503_ net599 vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__o21ai_1
X_05632_ net616 _01735_ _01736_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__or3_1
XANTENNA__08276__A core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06550__C1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08351_ _04431_ _04435_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05563_ net937 core.register_file.registers_state\[571\] net757 vssd1 vssd1 vccd1
+ vccd1 _01668_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07302_ _02967_ _02996_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08282_ _04374_ _04375_ net599 vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__o21ai_1
X_05494_ core.register_file.registers_state\[796\] core.register_file.registers_state\[828\]
+ core.register_file.registers_state\[924\] core.register_file.registers_state\[956\]
+ net707 net1019 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__05656__A1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07233_ core.register_file.registers_state\[289\] core.register_file.registers_state\[257\]
+ core.register_file.registers_state\[417\] core.register_file.registers_state\[385\]
+ net847 net1076 vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05839__S net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ _03267_ _03268_ net787 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06115_ net1046 core.register_file.registers_state\[840\] core.register_file.registers_state\[872\]
+ net677 net925 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__o221a_1
X_07095_ net767 _03187_ _03198_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o22a_4
XFILLER_0_100_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1037_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06046_ net935 core.register_file.registers_state\[74\] net693 core.register_file.registers_state\[106\]
+ net651 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout497_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout213 _04832_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout224 _04730_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
Xfanout235 _05248_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_4
XANTENNA__10165__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1204_A net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06908__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_4
XANTENNA__06908__B2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ net561 _04851_ net460 net272 net1686 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__a32o_1
Xfanout257 net260 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_6
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_8
X_07997_ net1113 _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout279 _05082_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06948_ _02242_ _02346_ _02521_ _02523_ _01632_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a41o_1
X_09736_ _04944_ net287 net274 net2163 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__a22o_1
XANTENNA__09858__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09322__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10523__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _04821_ net296 net284 net1967 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__a22o_1
X_06879_ _02981_ _02983_ net786 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout831_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06136__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07333__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08618_ _04673_ _04306_ _03964_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08186__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _04960_ net403 net301 net2013 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08617__C _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05895__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ core.pc.current_pc\[28\] core.pc.current_pc\[29\] _04603_ vssd1 vssd1 vccd1
+ vccd1 _04627_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11560_ clknet_leaf_26_clk _01072_ net1193 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05647__A1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511_ clknet_leaf_46_clk _00023_ net1290 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06844__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11491_ clknet_leaf_65_clk _01003_ net1245 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[963\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06705__Y _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10442_ net1389 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09389__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08125__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11029__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ net1450 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07495__S1 core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input58_A gpio_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11179__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09464__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 _01462_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_8
Xfanout791 _01455_ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__buf_4
XANTENNA__09849__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06168__X _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06532__C1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11827_ clknet_leaf_49_clk _01328_ net1310 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09616__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11758_ clknet_leaf_31_clk _00003_ net1205 vssd1 vssd1 vccd1 vccd1 core.ru.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08824__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06835__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10709_ clknet_leaf_62_clk _00221_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[181\]
+ sky130_fd_sc_hd__dfrtp_1
X_11689_ clknet_leaf_49_clk net1805 net1309 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06930__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload104 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06599__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07260__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07920_ net513 _03685_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nand2_2
XANTENNA__05810__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07851_ core.decoder.inst\[28\] net900 _03953_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10546__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ net1091 core.register_file.registers_state\[717\] core.register_file.registers_state\[749\]
+ net831 vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__o22a_1
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ _03762_ _03768_ net478 vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__mux2_2
XANTENNA__05407__B net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ _04822_ net401 net309 net2065 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a22o_1
XANTENNA__09304__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06733_ net813 _02836_ _02837_ net1088 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08718__B net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _04938_ net324 net314 net1971 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__a22o_1
X_06664_ net1109 core.register_file.registers_state\[212\] core.register_file.registers_state\[244\]
+ net859 net828 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__o221a_1
XFILLER_0_91_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08403_ _04492_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05615_ net938 core.register_file.registers_state\[951\] net757 net1010 vssd1 vssd1
+ vccd1 vccd1 _01720_ sky130_fd_sc_hd__o31a_1
X_09383_ net2093 net330 net323 _04806_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09068__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06595_ core.register_file.registers_state\[790\] core.register_file.registers_state\[822\]
+ net879 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ _02147_ _04430_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05546_ net1035 core.register_file.registers_state\[602\] vssd1 vssd1 vccd1 vccd1
+ _01651_ sky130_fd_sc_hd__or2_1
XANTENNA__06953__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08815__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08265_ _04354_ _04359_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05477_ net721 _01576_ _01581_ _01561_ _01567_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__o32a_4
XANTENNA_fanout412_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1154_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07216_ _01506_ _02451_ _02452_ net539 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ _01780_ _02718_ _03618_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05796__C net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07147_ core.register_file.registers_state\[548\] core.register_file.registers_state\[516\]
+ net854 vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08740__Y _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07784__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06054__A1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11321__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ core.register_file.registers_state\[806\] core.register_file.registers_state\[774\]
+ net841 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout781_A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08900__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06029_ net935 core.register_file.registers_state\[203\] net694 core.register_file.registers_state\[235\]
+ net636 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a221o_1
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_4
Xfanout1019 net1024 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_4
XANTENNA__10223__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__S0 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05317__B core.decoder.inst\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08909__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09719_ _04910_ net289 net274 net1937 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__a22o_1
X_10991_ clknet_leaf_82_clk _00503_ net1232 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06109__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05604__Y _01709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10310__A0 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07857__A2 _03959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05868__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05868__B2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11093__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11612_ clknet_leaf_27_clk _01124_ net1198 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08806__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07609__A2 _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11022__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08644__A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06817__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11543_ clknet_leaf_6_clk _01055_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1015\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06912__S0 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06293__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11474_ clknet_leaf_64_clk _00986_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[946\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10425_ net1356 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09231__A1 _04812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06045__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07242__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10356_ _05108_ net1597 net235 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__mux2_1
XANTENNA__09782__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10569__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10129__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10287_ net9 net902 net796 net2503 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05508__A _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06348__A2 _02451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06753__C1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09414__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05859__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05859__B2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05400_ net898 _01495_ _01503_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__nor3_4
XFILLER_0_5_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06380_ _02464_ _02471_ _02484_ net718 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__o22a_4
XANTENNA__08554__A _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05331_ core.ru.prev_busy core.ru.state\[3\] _01441_ vssd1 vssd1 vccd1 vccd1 _01444_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ net528 _04143_ _04154_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05262_ core.READ_I vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07001_ net807 _03104_ _03105_ net1085 vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__a211o_1
XANTENNA__05492__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10368__A0 _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06036__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09773__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__B1 _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ net2003 net369 _04941_ net437 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__a22o_1
XANTENNA__05795__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07540__A_N net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07903_ _03636_ _03707_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05418__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09525__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06013__S net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08883_ net243 net2394 net372 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
XANTENNA__10043__B net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _03635_ _03643_ _03653_ _03677_ net479 net496 vssd1 vssd1 vccd1 vccd1 _03939_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07765_ _03868_ _03869_ net482 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09504_ _04732_ net400 net309 net1791 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a22o_1
X_06716_ net793 _02817_ _02820_ net778 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07696_ _03645_ _03675_ net504 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__mux2_1
XANTENNA__06249__A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09435_ _04904_ net324 net314 net2099 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__a22o_1
X_06647_ _02750_ _02751_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_45_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1271_A net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout627_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09366_ net2010 net330 net324 _04707_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06578_ _02681_ _02682_ net1082 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08317_ net229 _04411_ _04412_ _04415_ _04360_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__o32a_1
X_05529_ net584 _01633_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__nor2_1
X_09297_ _04907_ net421 net334 net2039 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_X net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10071__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ core.pc.current_pc\[2\] _04352_ net598 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__mux2_1
XANTENNA__11598__Q core.IO_mod.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05483__C1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08179_ _03797_ _03959_ _03980_ _03950_ _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a221o_1
XANTENNA__10359__A0 _05111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08911__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ net1128 net2055 net913 _05213_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07224__B1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09764__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ clknet_leaf_61_clk _00702_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ _03862_ _05181_ net556 vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__a21o_1
XANTENNA__07527__B _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
Xoutput191 net191 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__09516__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ net1395 net517 _05142_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11274__RESET_B net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10974_ clknet_leaf_92_clk _00486_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07160__C1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__Y _04719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11367__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05710__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11526_ clknet_leaf_105_clk _01038_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[998\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_134_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05474__C1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ clknet_leaf_86_clk _00969_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[929\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07277__X _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10408_ net1329 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09409__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09755__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ clknet_leaf_42_clk _00900_ net1283 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[860\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ _02514_ net1502 net234 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__mux2_1
XANTENNA__10144__A _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09507__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07724__Y _03829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05880_ net629 _01983_ _01984_ net723 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_89_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07453__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07550_ net510 _03650_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08836__X _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09140__A0 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06501_ _02604_ _02605_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__nand2_1
XANTENNA__07377__S0 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07481_ net1104 core.register_file.registers_state\[863\] core.register_file.registers_state\[895\]
+ net850 net982 vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _04753_ net420 net341 net1708 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06432_ core.register_file.registers_state\[729\] core.register_file.registers_state\[761\]
+ net714 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09151_ _04910_ net351 net343 net1983 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06363_ core.register_file.registers_state\[290\] core.register_file.registers_state\[258\]
+ core.register_file.registers_state\[418\] core.register_file.registers_state\[386\]
+ net688 net1021 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08102_ net487 _03319_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__nor2_1
X_05314_ core.d_hit _01426_ _01423_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09082_ net2407 net366 net359 _04737_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06294_ net953 core.register_file.registers_state\[451\] vssd1 vssd1 vccd1 vccd1
+ _02399_ sky130_fd_sc_hd__and2_1
XANTENNA__09994__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ _04137_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput60 gpio_in[3] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xhold800 core.register_file.registers_state\[336\] vssd1 vssd1 vccd1 vccd1 net2119
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 core.ADR_I\[31\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout208_A _04334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06009__A1 _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07206__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 core.register_file.registers_state\[370\] vssd1 vssd1 vccd1 vccd1 net2141
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold833 core.register_file.registers_state\[50\] vssd1 vssd1 vccd1 vccd1 net2152
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold844 core.register_file.registers_state\[759\] vssd1 vssd1 vccd1 vccd1 net2163
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold855 core.register_file.registers_state\[721\] vssd1 vssd1 vccd1 vccd1 net2174
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold866 core.register_file.registers_state\[434\] vssd1 vssd1 vccd1 vccd1 net2185
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05419__Y _01524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 core.register_file.registers_state\[395\] vssd1 vssd1 vccd1 vccd1 net2196
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 core.register_file.registers_state\[421\] vssd1 vssd1 vccd1 vccd1 net2207
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ core.BUSY_O core.ru.state\[5\] net1129 vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold899 core.register_file.registers_state\[161\] vssd1 vssd1 vccd1 vccd1 net2218
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1117_A core.decoder.inst\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__C1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ net218 net735 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout577_A _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08866_ _04810_ net2449 net374 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__mux2_1
XANTENNA__08182__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07817_ _02519_ _03720_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nor2_2
X_08797_ core.IO_mod.input_reg\[25\] net251 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__and2_1
XANTENNA__06193__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07748_ _03660_ _03822_ net481 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08746__X _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A0 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout911_A _01449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07679_ net499 _03640_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__a21boi_1
XANTENNA__07142__C1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__B _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06496__A1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ net2341 _04815_ net405 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
X_10690_ clknet_leaf_78_clk _00202_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[162\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09349_ net1118 _04996_ net414 net1703 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__a22o_1
XANTENNA__06426__B _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09985__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout999_X net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ clknet_leaf_79_clk _00823_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09198__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ clknet_leaf_0_clk _00754_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[714\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09737__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11173_ clknet_leaf_100_clk _00685_ net1165 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[645\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input40_A gpio_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _03840_ _05170_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__and2_1
XANTENNA__11455__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ core.pc.current_pc\[2\] net591 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__or2_1
XANTENNA__10607__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09370__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09122__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05931__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ clknet_leaf_2_clk _00469_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[429\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05909__S1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07720__B net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10283__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08308__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10888_ clknet_leaf_13_clk _00400_ net1172 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[360\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05521__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08779__A3 _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08832__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ clknet_leaf_65_clk _01021_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[981\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_78_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold107 core.register_file.registers_state\[1018\] vssd1 vssd1 vccd1 vccd1 net1426
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 core.ADR_I\[24\] vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09189__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 core.ADR_I\[9\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09139__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09728__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07834__S1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08400__A2 _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 net610 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_2
XANTENNA__06411__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05845__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06981_ _03085_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_23_clk_X clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ net2060 net467 net433 _04782_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__a22o_1
X_05932_ net1054 core.register_file.registers_state\[142\] net681 core.register_file.registers_state\[174\]
+ net657 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_87_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10161__X _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11532__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1182 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09361__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08651_ _04717_ _04722_ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__and3_4
Xfanout1191 net1193 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_4
X_05863_ net964 _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__and2_1
XANTENNA__09900__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__C net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ net453 _02962_ net445 net503 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08582_ core.decoder.inst\[8\] net895 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_38_clk_X clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05794_ net1062 core.register_file.registers_state\[722\] core.register_file.registers_state\[754\]
+ net692 net662 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__o221a_1
XANTENNA__09113__A0 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07533_ _03636_ _03637_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07124__C1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06022__S0 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06478__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ core.register_file.registers_state\[31\] net678 net656 _03568_ vssd1 vssd1
+ vccd1 vccd1 _03569_ sky130_fd_sc_hd__a211o_1
XANTENNA__06527__A _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06415_ net554 _02381_ _02383_ net533 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__o211a_1
XANTENNA__05431__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09203_ _05010_ net361 net426 net1920 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09416__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07395_ core.register_file.registers_state\[793\] core.register_file.registers_state\[825\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1067_A core.decoder.inst\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ net205 core.register_file.registers_state\[215\] net347 vssd1 vssd1 vccd1
+ vccd1 _00255_ sky130_fd_sc_hd__mux2_1
XANTENNA__10026__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06346_ net720 _02434_ _02436_ _02444_ _02450_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__o32a_4
XANTENNA__08742__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ net742 net462 _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06277_ net586 _02347_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__nor2_2
XFILLER_0_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ net513 _03927_ _04017_ _04120_ _03688_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__o32a_1
XANTENNA__09719__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold630 core.register_file.registers_state\[560\] vssd1 vssd1 vccd1 vccd1 net1949
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 core.register_file.registers_state\[567\] vssd1 vssd1 vccd1 vccd1 net1960
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 core.register_file.registers_state\[500\] vssd1 vssd1 vccd1 vccd1 net1971
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold663 core.register_file.registers_state\[384\] vssd1 vssd1 vccd1 vccd1 net1982
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold674 core.register_file.registers_state\[889\] vssd1 vssd1 vccd1 vccd1 net1993
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold685 core.register_file.registers_state\[245\] vssd1 vssd1 vccd1 vccd1 net2004
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold696 core.register_file.registers_state\[506\] vssd1 vssd1 vccd1 vccd1 net2015
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05836__S0 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09967_ net1530 core.CPU_DAT_O\[23\] net801 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout861_A _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net563 _04918_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__and2_1
XANTENNA__09292__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ net1115 _05000_ net457 net378 net1527 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__a32o_1
XANTENNA__05606__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08849_ _04885_ net2322 net372 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__mux2_1
XANTENNA__10231__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11860_ clknet_leaf_28_clk net56 net1195 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08917__A _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10848__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10811_ clknet_leaf_19_clk _00323_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[283\]
+ sky130_fd_sc_hd__dfrtp_1
X_11791_ clknet_leaf_30_clk _01295_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06469__A1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10742_ clknet_leaf_44_clk _00254_ net1286 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[214\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10673_ clknet_leaf_75_clk _00185_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[145\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09407__A1 _04887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08652__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07969__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05487__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06641__A1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06172__A core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11225_ clknet_leaf_68_clk _00737_ net1267 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[697\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09591__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ clknet_leaf_57_clk _00668_ net1297 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[628\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ net471 _05162_ _05163_ net516 net1440 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__a32o_1
XANTENNA__05601__C1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ clknet_leaf_83_clk _00599_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[559\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05516__A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ net1595 net543 net522 _05119_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08697__A2 _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09894__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10589__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07106__C1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05380__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06004__S0 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06347__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05251__A core.decoder.inst\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06200_ core.register_file.registers_state\[518\] net674 net654 _02304_ vssd1 vssd1
+ vccd1 vccd1 _02305_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10008__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06880__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ _03281_ _03282_ _03284_ _03283_ net792 net827 vssd1 vssd1 vccd1 vccd1 _03285_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_76_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08082__A0 _03826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06131_ net1047 core.register_file.registers_state\[72\] core.register_file.registers_state\[104\]
+ net679 net641 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_65_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06093__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06632__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06062_ net1025 _02165_ _02166_ net1004 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a31o_1
XANTENNA__06632__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06082__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout406 net411 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_4
XANTENNA__09582__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_8
X_09821_ _04887_ net2377 net379 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
Xfanout428 net430 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_4
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10922__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09752_ _04973_ net289 net260 net1797 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__a22o_1
X_06964_ core.register_file.registers_state\[42\] core.register_file.registers_state\[10\]
+ net833 vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09334__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ core.IO_mod.input_reg\[10\] net253 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06021__S net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05915_ core.register_file.registers_state\[526\] net681 net658 _02019_ vssd1 vssd1
+ vccd1 vccd1 _02020_ sky130_fd_sc_hd__a211o_1
X_06895_ core.register_file.registers_state\[524\] core.register_file.registers_state\[556\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
XANTENNA__06148__B1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ net224 net2338 net280 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__mux2_1
XANTENNA__08688__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout275_A _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07896__B1 _03858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05846_ net960 _01950_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__nand2_1
X_08634_ net474 net544 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__and2_1
XANTENNA__08737__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08565_ net898 _01412_ core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__o21a_1
X_05777_ net1046 core.register_file.registers_state\[723\] core.register_file.registers_state\[755\]
+ net676 net652 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__o221a_1
XANTENNA__09637__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout442_A _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07516_ _01500_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__nor2_4
X_08496_ net228 _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ core.register_file.registers_state\[895\] net683 vssd1 vssd1 vccd1 vccd1
+ _03552_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06871__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07378_ net1108 core.register_file.registers_state\[345\] core.register_file.registers_state\[377\]
+ net858 net984 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06329_ _02427_ _02430_ net934 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__o21a_1
X_09117_ _04885_ net2364 net347 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11578__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06084__C1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ net613 net213 vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 core.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 core.register_file.registers_state\[804\] vssd1 vssd1 vccd1 vccd1 net1790
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08376__A1 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 core.register_file.registers_state\[400\] vssd1 vssd1 vccd1 vccd1 net1801
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ clknet_leaf_78_clk _00522_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07816__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09573__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold493 core.register_file.registers_state\[276\] vssd1 vssd1 vccd1 vccd1 net1812
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net941 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_2
XANTENNA__07535__B _02747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout951 net954 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout962 net963 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_4
XANTENNA__08128__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout973 _01371_ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08128__B2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09325__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06139__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 core.register_file.registers_state\[474\] vssd1 vssd1 vccd1 vccd1 net2479
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 core.register_file.registers_state\[177\] vssd1 vssd1 vccd1 vccd1 net2490
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 core.register_file.registers_state\[571\] vssd1 vssd1 vccd1 vccd1 net2501
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1193 core.register_file.registers_state\[130\] vssd1 vssd1 vccd1 vccd1 net2512
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07551__A _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11843_ clknet_leaf_36_clk net38 net1223 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05362__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09628__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07639__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08836__C1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ clknet_leaf_28_clk _01278_ net1194 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10725_ clknet_leaf_92_clk _00237_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[197\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06311__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07697__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10656_ clknet_leaf_53_clk _00168_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[128\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08064__A0 _03791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload16 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload16/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload27 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_6
X_10587_ clknet_leaf_19_clk _00099_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload38 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_12
XANTENNA__09800__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload49 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__inv_12
XANTENNA__06075__C1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07811__B1 _03915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06333__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09564__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09417__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ clknet_leaf_12_clk _00720_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ clknet_leaf_66_clk _00651_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[611\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08119__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07327__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05700_ _01798_ _01804_ net719 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a21o_1
X_06680_ _02782_ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07342__A2 _02534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire410_A _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05889__C1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05631_ net1040 core.register_file.registers_state\[215\] core.register_file.registers_state\[247\]
+ net671 net653 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__o221a_1
XANTENNA__06348__Y _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08350_ _04444_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05562_ net1040 net748 core.register_file.registers_state\[795\] vssd1 vssd1 vccd1
+ vccd1 _01667_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09095__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ _02999_ _03405_ _02966_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__o21ba_1
X_08281_ net209 _04381_ _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05493_ net633 _01595_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06302__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07232_ net967 _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07400__S net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ net995 core.register_file.registers_state\[195\] net885 core.register_file.registers_state\[227\]
+ net812 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06605__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06066__C1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06114_ net1007 _02213_ _02218_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06016__S net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ net776 _03192_ _03193_ net771 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__a31o_1
X_06045_ net637 _02149_ _02148_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_58_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09555__A0 _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout203 _04895_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
Xfanout214 _04820_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _04724_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
XANTENNA_fanout392_A _05066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 net240 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_4
Xfanout247 net248 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ net558 _04846_ net458 net270 net1722 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__a32o_1
XANTENNA__07030__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__B2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout258 net259 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10062__A _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout269 _05088_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_8
X_07996_ _02176_ _03081_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__or2_1
XANTENNA__11100__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _04942_ net296 net276 net1944 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__a22o_1
X_06947_ net771 _03045_ _03051_ _03040_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a31o_4
XANTENNA_fanout657_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ _04816_ net289 net282 net2382 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__a22o_1
X_06878_ core.register_file.registers_state\[14\] net877 net808 _02982_ vssd1 vssd1
+ vccd1 vccd1 _02983_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07371__A _03475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ _03884_ _03985_ _04004_ _04317_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__and4b_1
X_05829_ _01930_ _01931_ net622 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11250__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ _04959_ net399 net301 net2023 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__a22o_1
XANTENNA__08186__B _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_X net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08617__D _04317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ net228 _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__or2_1
XANTENNA__10818__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09086__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ core.pc.current_pc\[23\] _04558_ net231 vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08833__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08914__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ clknet_leaf_45_clk _00022_ net1289 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06844__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11490_ clknet_leaf_78_clk _01002_ net1253 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[962\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06715__A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10968__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ net1409 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09794__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10372_ net1468 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08061__A3 _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09745__B net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09546__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05765__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07546__A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 core.register_file.registers_state\[555\] vssd1 vssd1 vccd1 vccd1 net1609
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout770 _01469_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10863__RESET_B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout781 net783 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_8
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05583__A1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__A1 _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__A _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08521__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05353__X _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11826_ clknet_leaf_46_clk _01327_ net1290 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09700__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07088__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11757_ clknet_leaf_31_clk _00002_ net1201 vssd1 vssd1 vccd1 vccd1 core.ru.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06835__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ clknet_leaf_55_clk _00220_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[180\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11688_ clknet_leaf_32_clk _01200_ net1206 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06930__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload105 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__inv_6
X_10639_ clknet_leaf_82_clk _00151_ net1232 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09785__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07260__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06694__S0 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09537__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07012__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _01612_ _02660_ net580 _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__o211a_1
XANTENNA__07012__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06801_ _02875_ _02876_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06220__C1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07781_ _03812_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nand2_1
XANTENNA__11273__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
XANTENNA__10533__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09520_ _04817_ net397 net307 net1776 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__a22o_1
X_06732_ net996 core.register_file.registers_state\[690\] net887 core.register_file.registers_state\[658\]
+ net828 vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06663_ net1108 core.register_file.registers_state\[84\] core.register_file.registers_state\[116\]
+ net859 net813 vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__o221a_1
X_09451_ _04936_ net319 net312 net2487 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08402_ _01927_ _04491_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05614_ net938 core.register_file.registers_state\[823\] net757 net922 vssd1 vssd1
+ vccd1 vccd1 _01719_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09382_ net1771 net327 net317 _04801_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06594_ core.register_file.registers_state\[918\] core.register_file.registers_state\[950\]
+ net880 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
XANTENNA__09068__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08333_ core.pc.current_pc\[10\] _03080_ net576 vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05545_ net938 core.register_file.registers_state\[634\] net757 vssd1 vssd1 vccd1
+ vccd1 _01650_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08815__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10083__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08264_ _02347_ _04365_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_43_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06826__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05476_ net959 _01577_ _01580_ net628 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11392__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07215_ _03319_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__inv_2
X_08195_ _01781_ _02717_ net548 net900 net1019 vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__a32o_1
XANTENNA__11321__RESET_B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1147_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07146_ core.register_file.registers_state\[612\] core.register_file.registers_state\[580\]
+ net855 vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09776__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09240__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07251__A1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ core.register_file.registers_state\[934\] core.register_file.registers_state\[902\]
+ net839 vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09791__A3 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09528__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06028_ net935 core.register_file.registers_state\[75\] net693 core.register_file.registers_state\[107\]
+ net651 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_7_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_A _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1009 net1016 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07003__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07003__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05317__C net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _04080_ _04083_ net492 vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09718_ _04908_ net292 net277 net2086 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__a22o_1
XANTENNA__10640__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ clknet_leaf_88_clk _00502_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09700__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09649_ _04725_ net294 net285 net2157 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11611_ clknet_leaf_29_clk net1472 net1200 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10790__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08644__B _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06817__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11542_ clknet_leaf_61_clk _01054_ net1281 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1014\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08136__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06912__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11473_ clknet_leaf_90_clk _00985_ net1235 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[945\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07975__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09767__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ net1358 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08660__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09231__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07242__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10355_ _05107_ net1535 net233 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__mux2_1
XANTENNA__09519__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08990__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06450__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10129__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ net8 net903 net795 net2368 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__o22a_1
XANTENNA__06180__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05508__B _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05556__A1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05524__A _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08835__A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09430__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ clknet_leaf_54_clk _01310_ net1299 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_107_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08554__B _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05330_ core.ru.prev_busy _01441_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05261_ net1013 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XANTENNA__06284__A2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07481__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07481__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07000_ net997 core.register_file.registers_state\[681\] net872 core.register_file.registers_state\[649\]
+ net821 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09758__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__X _03843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09222__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10513__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06667__S0 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09773__A3 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10785__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08981__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ net573 _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06992__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07902_ _02968_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_36_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05418__B net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08882_ net203 net2469 net371 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11789__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09930__A0 core.decoder.inst\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07833_ net511 _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_32_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07764_ _03803_ _03805_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09503_ _04726_ net400 net309 net1685 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06715_ net788 _02818_ _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__or3_1
X_07695_ net497 _03671_ _03799_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ _04902_ net323 net314 net2251 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06646_ _02747_ _02749_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__nand2_1
XANTENNA__06964__S net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09365_ net566 _05030_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout522_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06577_ net1095 core.register_file.registers_state\[471\] core.register_file.registers_state\[503\]
+ net836 net1071 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ _04413_ _04414_ net597 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05528_ core.decoder.inst\[26\] net898 net593 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ _04905_ net421 net334 net2150 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__a22o_1
XANTENNA__09461__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08247_ _04351_ _01380_ net230 vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07472__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05459_ net653 _01554_ _01563_ net1005 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07472__B2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_X net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08178_ _03773_ _03949_ _04280_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout891_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08016__A3 _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__A2 _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout989_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ _03231_ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__and2_1
XANTENNA__06658__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10140_ _03862_ _05181_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__nor2_1
XANTENNA__07096__A _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05786__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XANTENNA__07527__C net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput192 net192 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_10071_ _04139_ net557 net590 core.pc.current_pc\[8\] net472 vssd1 vssd1 vccd1 vccd1
+ _05142_ sky130_fd_sc_hd__o221a_1
XANTENNA__05328__B core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09921__A0 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05538__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05538__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__B _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10973_ clknet_leaf_19_clk _00485_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[445\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07160__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05710__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05350__Y _01455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06175__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__X _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09452__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ clknet_leaf_86_clk _01037_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[997\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_135_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06671__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ clknet_leaf_57_clk _00968_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[928\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09204__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10407_ net1334 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11387_ clknet_leaf_23_clk _00899_ net1184 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10338_ _02451_ net1491 net234 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
XANTENNA__05777__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06974__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05777__B2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10269_ core.BUSY_O wb.prev_BUSY_O net902 vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and3b_1
XANTENNA__09425__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05254__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08479__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06500_ _01488_ _02603_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__nand2_1
XANTENNA__10286__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07377__S1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07480_ net1104 core.register_file.registers_state\[991\] core.register_file.registers_state\[1023\]
+ net850 net1077 vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05541__X _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06431_ core.register_file.registers_state\[665\] core.register_file.registers_state\[697\]
+ net712 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10038__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05260__Y _01375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06362_ net1059 core.register_file.registers_state\[482\] net755 _02466_ vssd1 vssd1
+ vccd1 vccd1 _02467_ sky130_fd_sc_hd__a31o_1
X_09150_ _04908_ net357 net345 net2173 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09443__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05313_ core.d_hit _01426_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08101_ net1113 _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11461__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06293_ net1060 core.register_file.registers_state\[355\] net754 _02397_ vssd1 vssd1
+ vccd1 vccd1 _02398_ sky130_fd_sc_hd__a31o_1
X_09081_ net2328 net366 net359 _04731_ vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ net506 _03701_ _03752_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput50 gpio_in[23] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput61 gpio_in[4] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08504__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold801 core.register_file.registers_state\[188\] vssd1 vssd1 vccd1 vccd1 net2120
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold812 core.register_file.registers_state\[321\] vssd1 vssd1 vccd1 vccd1 net2131
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07206__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold823 core.register_file.registers_state\[463\] vssd1 vssd1 vccd1 vccd1 net2142
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold834 core.register_file.registers_state\[858\] vssd1 vssd1 vccd1 vccd1 net2153
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold845 core.register_file.registers_state\[641\] vssd1 vssd1 vccd1 vccd1 net2164
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold856 core.register_file.registers_state\[334\] vssd1 vssd1 vccd1 vccd1 net2175
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 core.register_file.registers_state\[489\] vssd1 vssd1 vccd1 vccd1 net2186
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold878 core.register_file.registers_state\[815\] vssd1 vssd1 vccd1 vccd1 net2197
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ core.ru.state\[0\] core.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__nor2_1
Xhold889 core.register_file.registers_state\[354\] vssd1 vssd1 vccd1 vccd1 net2208
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05768__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05768__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06251__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08934_ net2260 net369 _04929_ net436 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1012_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08865_ _04805_ net2494 net374 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout472_A _05127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07816_ net512 _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__nor2_1
XANTENNA__06193__A1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08796_ net1882 net466 net435 _04846_ vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__a22o_1
XANTENNA__11754__RESET_B net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ core.decoder.inst\[29\] net899 _03849_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_
+ sky130_fd_sc_hd__a211o_2
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10277__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07678_ net455 _02717_ net447 net497 vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08906__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ core.register_file.registers_state\[466\] net216 net408 vssd1 vssd1 vccd1
+ vccd1 _00506_ sky130_fd_sc_hd__mux2_1
XANTENNA__06496__A2 _01709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06629_ net1105 core.register_file.registers_state\[181\] net851 core.register_file.registers_state\[149\]
+ net810 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1267_X net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09348_ net1115 _04994_ net412 net1801 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09434__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10229__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ net2345 _04815_ net335 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
XANTENNA__05456__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11310_ clknet_leaf_81_clk _00822_ net1235 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[782\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07819__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06653__C1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08414__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05551__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ clknet_leaf_17_clk _00753_ net1211 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[713\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06405__C1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11522__SET_B net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ clknet_leaf_80_clk _00684_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[644\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10123_ _03840_ _05170_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10054_ net471 _05130_ _05131_ net516 net1613 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__a32o_1
XANTENNA__07554__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__S0 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05931__A1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10956_ clknet_leaf_102_clk _00468_ net1162 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[428\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09673__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07684__A1 _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10887_ clknet_leaf_93_clk _00399_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[359\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07436__A1 _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08633__B1 _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__B net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07987__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ clknet_leaf_51_clk _01020_ net1297 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[980\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05998__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05998__B2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 core.register_file.registers_state\[974\] vssd1 vssd1 vccd1 vccd1 net1427
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 core.register_file.registers_state\[14\] vssd1 vssd1 vccd1 vccd1 net1438
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ clknet_leaf_83_clk _00951_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10155__A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06411__A2 _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06980_ _03083_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__and2_1
XANTENNA__05845__S1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05931_ net964 _02022_ _02027_ net718 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_87_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05255__Y _01370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1170 net1171 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
X_08650_ net728 _04215_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__nand2_1
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_2
Xfanout1192 net1193 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
X_05862_ core.register_file.registers_state\[273\] core.register_file.registers_state\[305\]
+ core.register_file.registers_state\[401\] core.register_file.registers_state\[433\]
+ net711 net1020 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__mux4_1
X_07601_ net453 _02994_ net445 net508 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__a31o_1
XANTENNA__07751__X _03856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08581_ core.decoder.inst\[7\] net895 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__nand2_2
XANTENNA__05922__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05793_ net1062 core.register_file.registers_state\[594\] core.register_file.registers_state\[626\]
+ net692 net648 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__o221a_1
X_07532_ net452 _02873_ net444 net502 vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09664__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05712__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06022__S1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07463_ net1053 core.register_file.registers_state\[63\] net751 vssd1 vssd1 vccd1
+ vccd1 _03568_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09202_ _05008_ net353 net423 net1635 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__a22o_1
X_06414_ net493 net476 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10851__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06019__S net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07394_ _03495_ _03496_ _03497_ _03498_ net793 net813 vssd1 vssd1 vccd1 vccd1 _03499_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10049__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09133_ net213 net2061 net349 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07427__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06345_ net634 _02446_ _02449_ net723 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07427__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08742__B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06276_ _02372_ _02379_ _02364_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a21o_1
X_09064_ net613 net210 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08015_ _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__inv_2
XANTENNA__10065__A _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold620 net168 vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 core.register_file.registers_state\[234\] vssd1 vssd1 vccd1 vccd1 net1950
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold642 core.register_file.registers_state\[729\] vssd1 vssd1 vccd1 vccd1 net1961
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold653 core.register_file.registers_state\[885\] vssd1 vssd1 vccd1 vccd1 net1972
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 core.register_file.registers_state\[230\] vssd1 vssd1 vccd1 vccd1 net1983
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 core.register_file.registers_state\[678\] vssd1 vssd1 vccd1 vccd1 net1994
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 core.register_file.registers_state\[143\] vssd1 vssd1 vccd1 vccd1 net2005
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout687_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 core.register_file.registers_state\[382\] vssd1 vssd1 vccd1 vccd1 net2016
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ net1494 core.CPU_DAT_O\[22\] net800 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__mux2_1
XANTENNA__05836__S1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06689__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1015_X net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07374__A _03475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08917_ _04769_ net601 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__nor2_1
X_09897_ net1119 _05075_ net376 net1696 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__a22o_1
XANTENNA__08189__B _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09352__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05606__B _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ _04656_ _04746_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06166__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08779_ net728 _04830_ _04831_ _04829_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__o31a_2
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05374__C1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08917__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10810_ clknet_leaf_9_clk _00322_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[282\]
+ sky130_fd_sc_hd__dfrtp_1
X_11790_ clknet_leaf_29_clk _01294_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07115__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09655__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08863__A0 _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ clknet_leaf_64_clk _00253_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[213\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05677__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10888__RESET_B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10672_ clknet_leaf_108_clk _00184_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[144\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08933__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08652__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05429__B1 _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06172__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07983__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11224_ clknet_leaf_3_clk _00736_ net1150 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06929__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07051__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ clknet_leaf_11_clk _00667_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[627\]
+ sky130_fd_sc_hd__dfrtp_1
X_10106_ _04306_ net589 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__nand2_1
XANTENNA_input36_X net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ clknet_leaf_82_clk _00598_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[558\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09343__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
X_10037_ net594 _01582_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__nor2_1
XANTENNA__08667__X _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09004__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05532__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06004__S1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10256__A3 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ clknet_leaf_19_clk _00451_ net1191 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[411\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06347__B _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06865__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10558__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
X_06130_ net656 _02233_ _02234_ net617 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__o211a_1
XANTENNA__06617__C1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08082__A1 _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06061_ net935 core.register_file.registers_state\[714\] net693 core.register_file.registers_state\[746\]
+ net636 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _04886_ net2272 net380 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
Xfanout407 net410 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_6
Xfanout418 _05029_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_6
XANTENNA__10192__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _04971_ net292 net259 net1942 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__a22o_1
XANTENNA__05707__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06963_ net1093 core.register_file.registers_state\[138\] net833 core.register_file.registers_state\[170\]
+ net817 vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_78_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_08702_ core.IO_mod.data_from_mem\[10\] net247 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__nand2_1
XANTENNA__09334__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05914_ net1054 core.register_file.registers_state\[558\] net753 vssd1 vssd1 vccd1
+ vccd1 _02019_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ net225 net2337 net280 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__mux2_1
XANTENNA__06148__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06894_ _02966_ _02967_ _02998_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__or3_1
XANTENNA__09885__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ core.decoder.inst\[11\] _04661_ _04662_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_96_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05845_ core.register_file.registers_state\[272\] core.register_file.registers_state\[304\]
+ core.register_file.registers_state\[400\] core.register_file.registers_state\[432\]
+ net695 net1013 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08564_ core.pc.current_pc\[30\] net595 _04638_ _04640_ vssd1 vssd1 vccd1 vccd1 _00038_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09098__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05776_ net627 _01875_ net722 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07133__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07515_ _01400_ _01619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__or2_2
XANTENNA__08845__A0 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ _04556_ _04575_ _04574_ _04565_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_18_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout435_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05659__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07446_ core.register_file.registers_state\[1023\] net683 vssd1 vssd1 vccd1 vccd1
+ _03551_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout602_A _04897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout223_X net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ core.register_file.registers_state\[281\] core.register_file.registers_state\[313\]
+ core.register_file.registers_state\[409\] core.register_file.registers_state\[441\]
+ net889 net1080 vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06608__C1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ _04884_ net2227 net349 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06328_ net955 core.register_file.registers_state\[832\] net713 core.register_file.registers_state\[864\]
+ net1022 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09047_ net2360 net429 _05004_ net437 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__a22o_1
X_06259_ net634 _02363_ _02358_ net718 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a211oi_1
XANTENNA__10304__A_N _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05831__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold450 core.register_file.registers_state\[445\] vssd1 vssd1 vccd1 vccd1 net1769
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout971_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 core.register_file.registers_state\[821\] vssd1 vssd1 vccd1 vccd1 net1780
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold472 core.register_file.registers_state\[547\] vssd1 vssd1 vccd1 vccd1 net1791
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold483 core.register_file.registers_state\[418\] vssd1 vssd1 vccd1 vccd1 net1802
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07816__B _03920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold494 core.register_file.registers_state\[924\] vssd1 vssd1 vccd1 vccd1 net1813
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10183__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_2
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_4
X_09949_ core.IO_mod.data_from_mem\[5\] net2483 net798 vssd1 vssd1 vccd1 vccd1 _01101_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout952 net953 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_2
XANTENNA__07535__C net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout963 net966 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__buf_4
XFILLER_0_95_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08128__A2 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout974 net975 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_4
Xfanout985 _01370_ vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_4
Xhold1150 core.register_file.registers_state\[93\] vssd1 vssd1 vccd1 vccd1 net2469
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09876__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1161 core.register_file.registers_state\[265\] vssd1 vssd1 vccd1 vccd1 net2480
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 core.register_file.registers_state\[845\] vssd1 vssd1 vccd1 vccd1 net2491
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 core.register_file.registers_state\[210\] vssd1 vssd1 vccd1 vccd1 net2502
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 core.register_file.registers_state\[720\] vssd1 vssd1 vccd1 vccd1 net2513
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05898__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11842_ clknet_leaf_35_clk net37 net1208 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08139__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__A3 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ clknet_leaf_24_clk _01277_ net1184 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07978__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10724_ clknet_leaf_77_clk _00236_ net1261 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[196\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06311__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_22_clk_X clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ clknet_leaf_94_clk _00167_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload17 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_114_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload28 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_6
X_10586_ clknet_leaf_9_clk _00098_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09800__A2 _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload39 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__07811__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05822__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11672__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ clknet_leaf_91_clk _00719_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[679\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07024__C1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10174__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__B1 core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11138_ clknet_leaf_80_clk _00650_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[610\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06122__S net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ clknet_leaf_17_clk _00581_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[541\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_0_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09867__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07878__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05630_ net1039 core.register_file.registers_state\[87\] core.register_file.registers_state\[119\]
+ net671 net638 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06550__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06358__A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06550__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05984__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05561_ net1040 net748 core.register_file.registers_state\[923\] vssd1 vssd1 vccd1
+ vccd1 _01666_ sky130_fd_sc_hd__a21o_1
XANTENNA__08827__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07300_ _02935_ _03404_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08280_ _04376_ _04378_ _04379_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__or3_1
X_05492_ net962 _01586_ _01596_ net628 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06302__A1 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07231_ net1086 _03334_ _03335_ _03333_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07162_ net995 core.register_file.registers_state\[67\] net885 core.register_file.registers_state\[99\]
+ net827 vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06113_ _02215_ _02216_ _02217_ _02214_ net932 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07263__C1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07093_ net1084 _03194_ _03197_ net780 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05813__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06044_ core.register_file.registers_state\[42\] core.register_file.registers_state\[10\]
+ net668 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06380__X _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07015__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout204 _04894_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout215 _04815_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
XANTENNA__10165__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09803_ net559 _04840_ net456 net270 net2075 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__a32o_1
Xfanout237 net240 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_2
XANTENNA__10062__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ _04078_ _04081_ _04082_ _04099_ net494 net481 vssd1 vssd1 vccd1 vccd1 _04100_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_66_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout385_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__Y _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _04940_ net296 net276 net2135 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__a22o_1
XANTENNA__07688__A2_N net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06946_ net1083 _03049_ _03050_ net1066 _03048_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a311o_1
XFILLER_0_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09858__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ _04811_ net296 net284 net2274 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__a22o_1
X_06877_ core.register_file.registers_state\[46\] net847 vssd1 vssd1 vccd1 vccd1 _02982_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ net732 net253 core.IO_mod.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 _04691_
+ sky130_fd_sc_hd__a21o_2
X_05828_ core.register_file.registers_state\[528\] core.register_file.registers_state\[560\]
+ net697 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
X_09596_ _04957_ net396 net299 net2139 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08547_ _04620_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__xor2_1
XANTENNA__08818__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05759_ _01862_ _01863_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_X net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07798__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ core.pc.current_pc\[22\] core.pc.current_pc\[23\] _04540_ vssd1 vssd1 vccd1
+ vccd1 _04562_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09491__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07429_ net970 _03530_ _03533_ net775 vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05501__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__A _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10440_ net1347 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09243__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10237__B net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07254__C1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ net1439 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08930__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08422__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout974_X net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 core.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10253__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold291 core.register_file.registers_state\[388\] vssd1 vssd1 vccd1 vccd1 net1610
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10156__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 net762 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_4
Xfanout771 _01468_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_8
Xfanout782 net783 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout793 net794 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09849__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06178__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11825_ clknet_leaf_70_clk _01326_ net1274 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08809__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11756_ clknet_leaf_31_clk _00001_ net1205 vssd1 vssd1 vccd1 vccd1 core.ru.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_79_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06296__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ clknet_leaf_97_clk _00219_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[179\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10912__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ clknet_leaf_49_clk _01199_ net1310 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09001__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10638_ clknet_leaf_90_clk _00150_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09234__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload106 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__inv_12
XFILLER_0_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06048__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10569_ clknet_leaf_40_clk _00081_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06599__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09428__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06694__S1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05257__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ _02848_ _02903_ _02904_ _02814_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__o211a_2
XANTENNA__06220__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07780_ _03421_ _03422_ _03540_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_1
X_06731_ core.register_file.registers_state\[530\] core.register_file.registers_state\[562\]
+ net887 vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09450_ _04934_ net324 net313 net2417 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a22o_1
X_06662_ core.register_file.registers_state\[20\] core.register_file.registers_state\[52\]
+ net890 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__mux2_1
XANTENNA__06523__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ _01927_ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05613_ net642 _01714_ _01715_ _01716_ _01717_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a32o_1
X_09381_ net1807 net329 net322 _04796_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06593_ core.register_file.registers_state\[982\] core.register_file.registers_state\[1014\]
+ net880 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08332_ _04427_ _04428_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05544_ net939 core.register_file.registers_state\[698\] net696 core.register_file.registers_state\[666\]
+ net653 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09473__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07411__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06287__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08263_ _02347_ _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_43_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07484__C1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05475_ _01578_ _01579_ net1026 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07214_ net774 _03318_ _03305_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__o21a_4
XFILLER_0_7_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08194_ _03413_ _03416_ _03419_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__nor3_1
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09225__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06039__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07145_ core.register_file.registers_state\[740\] core.register_file.registers_state\[708\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07076_ _03177_ _03178_ _03179_ _03180_ net790 net819 vssd1 vssd1 vccd1 vccd1 _03181_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_7_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09528__A1 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06027_ _02129_ _02131_ net616 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_7_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1307_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08200__A1 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11098__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ _04081_ _04082_ net485 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux2_1
XANTENNA__05317__D net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05565__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ _04906_ net294 net276 net1931 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__a22o_1
X_06929_ net789 _03032_ _03033_ net779 vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout934_A _01375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09648_ _04720_ net292 net284 net2103 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__a22o_1
XANTENNA__08765__X _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08621__D_N _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07711__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _04923_ net397 net299 net1859 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__a22o_1
X_11610_ clknet_leaf_33_clk _01122_ net1204 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06726__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11541_ clknet_leaf_65_clk _01053_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1013\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07475__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ clknet_leaf_103_clk _00984_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[944\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09216__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06293__A3 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__C1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ net1333 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08660__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input63_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _05106_ net1515 net232 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__mux2_1
XANTENNA__06461__A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09519__A1 _04812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08990__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10285_ net7 net904 net797 core.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_109_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06753__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net592 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_2
XANTENNA__06753__B2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09711__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08835__B net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11808_ clknet_leaf_49_clk _01309_ net1309 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09455__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09012__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11739_ clknet_leaf_37_clk _01251_ net1222 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07466__C1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05260_ net1005 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkinv_4
XANTENNA__09207__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05492__A1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06642__Y _02747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06036__A3 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08430__A1 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__S1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05258__Y _01373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ _04826_ net602 vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__nor2_2
XANTENNA__06992__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10808__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ _02935_ _02998_ _04005_ _02996_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__o31a_1
XFILLER_0_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08881_ net741 _04870_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07832_ _03638_ _03708_ _03711_ _03700_ net485 net490 vssd1 vssd1 vccd1 vccd1 _03937_
+ sky130_fd_sc_hd__mux4_2
X_07763_ net497 _03671_ _03806_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__o21a_1
XANTENNA__05952__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ net569 _04720_ net399 net310 net1620 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06714_ net1108 core.register_file.registers_state\[210\] core.register_file.registers_state\[242\]
+ net858 net829 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__o221a_1
XANTENNA__09694__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07694_ net451 _03506_ net443 net504 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ _04900_ net321 net313 net2101 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__a22o_1
XANTENNA__06249__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06645_ _02747_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__nor2_1
XANTENNA__05704__C1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__A1 _03289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _05022_ _05030_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__or2_4
XANTENNA__09446__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06576_ net1095 core.register_file.registers_state\[343\] core.register_file.registers_state\[375\]
+ net836 net979 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08315_ core.pc.current_pc\[8\] _04403_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__nor2_1
X_05527_ net581 _01630_ _01628_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__or3b_4
X_09295_ _04903_ net421 net334 net2208 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout515_A _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1257_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _04341_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05458_ net942 core.register_file.registers_state\[701\] net762 vssd1 vssd1 vccd1
+ vccd1 _01563_ sky130_fd_sc_hd__or3_1
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08761__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05483__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07209__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08177_ net1112 _01864_ net551 _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__o31a_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05389_ _01493_ _01392_ _01400_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__A3 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ _02346_ _03232_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06658__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout884_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07059_ net1088 _03162_ _03163_ net967 vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a31o_1
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__clkbuf_4
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_101_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_10070_ net1552 net518 _05141_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__a21o_1
Xoutput193 net193 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06196__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05943__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10972_ clknet_leaf_40_clk _00484_ net1216 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[444\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08936__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10295__A1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05912__X _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07160__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11113__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09988__B2 _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11524_ clknet_leaf_81_clk _01036_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[996\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_68_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire221 _04790_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
XFILLER_0_110_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05474__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11283__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05474__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11455_ clknet_leaf_15_clk _00967_ net1177 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[927\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ net1331 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11386_ clknet_leaf_6_clk _00898_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ _04229_ net245 vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__nand2_4
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06974__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07574__X _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10268_ wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__nand2_1
XANTENNA__08176__B1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ net79 net914 vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_128_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07226__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09007__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06918__X _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08846__A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06430_ core.decoder.inst\[25\] net899 net593 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06361_ net952 core.register_file.registers_state\[450\] vssd1 vssd1 vccd1 vccd1
+ _02466_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08852__Y _04887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ net487 _03319_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05312_ _01406_ _01417_ _01425_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__or3_4
X_09080_ net2435 net366 net359 _04725_ vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__a22o_1
X_06292_ net953 core.register_file.registers_state\[323\] net1020 vssd1 vssd1 vccd1
+ vccd1 _02397_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08581__A core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08031_ _03658_ _03891_ _04129_ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__o211a_1
Xinput40 gpio_in[14] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
Xhold802 core.register_file.registers_state\[457\] vssd1 vssd1 vccd1 vccd1 net2121
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10630__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold813 core.register_file.registers_state\[672\] vssd1 vssd1 vccd1 vccd1 net2132
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09600__A0 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold824 core.register_file.registers_state\[738\] vssd1 vssd1 vccd1 vccd1 net2143
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold835 core.register_file.registers_state\[648\] vssd1 vssd1 vccd1 vccd1 net2154
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold846 core.register_file.registers_state\[135\] vssd1 vssd1 vccd1 vccd1 net2165
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold857 core.register_file.registers_state\[173\] vssd1 vssd1 vccd1 vccd1 net2176
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09982_ net727 _01426_ core.d_hit _01367_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a211oi_4
Xhold868 core.register_file.registers_state\[341\] vssd1 vssd1 vccd1 vccd1 net2187
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold879 core.register_file.registers_state\[745\] vssd1 vssd1 vccd1 vccd1 net2198
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ net572 net219 net737 vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_A _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ net218 net2406 net371 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1005_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ _03704_ _03724_ _03728_ _03717_ net483 net490 vssd1 vssd1 vccd1 vccd1 _03920_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_93_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05925__C1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ net564 net606 _04844_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07746_ net1114 _03848_ _03850_ net580 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__o211a_1
XANTENNA__08014__S0 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_A _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07142__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ net2350 net217 net408 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06628_ net777 _02731_ _02732_ net773 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__o211a_1
X_09347_ net1119 _04992_ net414 net1630 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06559_ net1094 core.register_file.registers_state\[855\] core.register_file.registers_state\[887\]
+ net835 net979 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ net2369 net216 net337 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ net228 vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05551__S1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ clknet_leaf_13_clk _00752_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09198__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10245__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06405__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11171_ clknet_leaf_66_clk _00683_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[643\]
+ sky130_fd_sc_hd__dfrtp_1
X_10122_ net470 _05171_ _05174_ net515 net1435 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10053_ _04229_ net589 vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__nand2_1
XANTENNA__07554__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__S1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05916__C1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07381__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09658__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09261__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10503__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955_ clknet_leaf_108_clk _00467_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[427\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07684__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10886_ clknet_leaf_105_clk _00398_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[358\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10653__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07436__A2 _03422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09830__A0 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08633__A1 core.decoder.inst\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ clknet_leaf_11_clk _01019_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[979\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08832__C net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__B _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09189__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 core.register_file.registers_state\[1016\] vssd1 vssd1 vccd1 vccd1 net1428
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11438_ clknet_leaf_81_clk _00950_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11369_ clknet_leaf_38_clk _00881_ net1213 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[841\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06947__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05964__S net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__A _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05930_ _02030_ _02034_ net964 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11159__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09897__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1167 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_4
Xfanout1171 net1172 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09361__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05861_ _01962_ _01965_ net634 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a21o_1
Xfanout1182 net1209 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__buf_2
XANTENNA__05907__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1209 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_2
X_07600_ _03700_ _03704_ net486 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__mux2_1
X_08580_ core.decoder.inst\[7\] net895 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and2_4
X_05792_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__inv_2
XANTENNA__09649__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08576__A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06580__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire221_X net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ net452 _02900_ net444 net508 vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07124__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07462_ net1053 core.register_file.registers_state\[191\] net678 core.register_file.registers_state\[159\]
+ net641 vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_27_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08600__A_N _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06332__C1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ net603 net205 net352 net423 net1749 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__a32o_1
X_06413_ net487 net482 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__nor2_2
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05431__C net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07393_ core.register_file.registers_state\[601\] core.register_file.registers_state\[633\]
+ net888 vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11134__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ _04891_ net2031 net349 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__mux2_1
X_06344_ _02447_ _02448_ net965 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08624__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__A0 _04887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09063_ net2231 net427 _05014_ net432 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06275_ _02372_ _02379_ _02364_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout213_A _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08014_ _04008_ _04055_ _04057_ _04117_ net496 net480 vssd1 vssd1 vccd1 vccd1 _04119_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_103_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold610 core.register_file.registers_state\[530\] vssd1 vssd1 vccd1 vccd1 net1929
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold621 core.register_file.registers_state\[365\] vssd1 vssd1 vccd1 vccd1 net1940
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10065__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold632 core.register_file.registers_state\[891\] vssd1 vssd1 vccd1 vccd1 net1951
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 core.register_file.registers_state\[708\] vssd1 vssd1 vccd1 vccd1 net1962
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold654 core.register_file.registers_state\[766\] vssd1 vssd1 vccd1 vccd1 net1973
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10195__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 core.register_file.registers_state\[795\] vssd1 vssd1 vccd1 vccd1 net1984
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06399__C1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 core.register_file.registers_state\[865\] vssd1 vssd1 vccd1 vccd1 net1995
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05874__S net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 core.register_file.registers_state\[52\] vssd1 vssd1 vccd1 vccd1 net2006
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 core.register_file.registers_state\[123\] vssd1 vssd1 vccd1 vccd1 net2017
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ net2209 core.CPU_DAT_O\[21\] net801 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout582_A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net2346 net368 _04917_ net434 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__a22o_1
X_09896_ net1119 _05074_ net376 net1702 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__a22o_1
XANTENNA__09888__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_X net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10526__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ _04884_ net2247 net373 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ core.IO_mod.data_from_mem\[22\] net248 vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06571__C1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ net510 _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10740_ clknet_leaf_53_clk _00252_ net1302 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[212\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10676__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06323__C1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05677__A1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10671_ clknet_leaf_84_clk _00183_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[143\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08933__B net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08076__C1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11223_ clknet_leaf_9_clk _00735_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[695\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07836__Y _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10186__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06929__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11301__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07051__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09591__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ clknet_leaf_68_clk _00666_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[626\]
+ sky130_fd_sc_hd__dfrtp_1
X_10105_ core.pc.current_pc\[22\] net589 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__or2_1
XANTENNA__05601__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__A0 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11085_ clknet_leaf_2_clk _00597_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[557\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10036_ net1499 net543 net522 _05118_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__a22o_1
XANTENNA__11451__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05460__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07106__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07106__B2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09004__B _04975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10938_ clknet_leaf_8_clk _00450_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[410\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06865__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10869_ clknet_leaf_61_clk _00381_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[341\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06644__A _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06712__S0 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06093__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06060_ net935 core.register_file.registers_state\[586\] net693 core.register_file.registers_state\[618\]
+ net651 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05840__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10177__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire550_A _02810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout408 net409 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_4
XANTENNA__09582__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A2_N _04018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout419 net420 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
XANTENNA__08790__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _04969_ net294 net258 net1867 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__a22o_1
X_06962_ _03061_ _03066_ net779 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
X_08701_ net732 _04109_ net526 vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__o21ai_1
X_05913_ net585 _02017_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__nor2_1
X_09681_ net226 net2256 net281 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06893_ _02996_ _02997_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08632_ net608 net207 vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__and2_2
X_05844_ net621 _01945_ _01948_ net628 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07414__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08737__C _04795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ net208 _04639_ net595 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__o21ai_1
X_05775_ net960 _01876_ _01879_ net627 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a211o_1
XANTENNA__11315__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ net898 net580 vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _04574_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__nor2_1
XANTENNA__07648__A2 _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06305__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__X _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ _02635_ _02662_ _03548_ _02633_ _02606_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__a311o_2
XFILLER_0_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout330_A _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout428_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ _03451_ _03480_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09115_ _04736_ net2456 net350 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06327_ net955 core.register_file.registers_state\[960\] net713 core.register_file.registers_state\[992\]
+ net930 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06084__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09046_ net573 _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06258_ _02359_ _02360_ _02361_ _02362_ net623 net660 vssd1 vssd1 vccd1 vccd1 _02363_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05831__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 net155 vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ net1027 _02291_ _02293_ net627 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10168__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1125_X net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 net192 vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 core.register_file.registers_state\[522\] vssd1 vssd1 vccd1 vccd1 net1781
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 core.register_file.registers_state\[890\] vssd1 vssd1 vccd1 vccd1 net1792
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 core.register_file.registers_state\[527\] vssd1 vssd1 vccd1 vccd1 net1803
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold495 core.register_file.registers_state\[623\] vssd1 vssd1 vccd1 vccd1 net1814
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_2
Xfanout931 _01376_ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__buf_4
X_09948_ net2116 core.CPU_DAT_O\[4\] net800 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
Xfanout942 net943 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_2
XANTENNA__06792__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout975 _01371_ vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_4
XANTENNA__09325__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_2
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _04704_ net2127 net376 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__mux2_1
Xfanout997 _01369_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__buf_6
XANTENNA__06139__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1140 core.register_file.registers_state\[603\] vssd1 vssd1 vccd1 vccd1 net2459
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 core.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 core.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05347__B1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 core.register_file.registers_state\[217\] vssd1 vssd1 vccd1 vccd1 net2492
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10340__A0 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06544__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1184 core.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_120_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05898__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1195 core.register_file.registers_state\[350\] vssd1 vssd1 vccd1 vccd1 net2514
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11841_ clknet_leaf_35_clk net36 net1220 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09628__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09599__X _05066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07639__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11772_ clknet_leaf_24_clk _01276_ net1187 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08944__A _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10723_ clknet_leaf_71_clk _00235_ net1270 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[195\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06735__Y _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10654_ clknet_leaf_96_clk _00166_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09261__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ clknet_leaf_69_clk _00097_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload18 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload18/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__08950__Y _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload29 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_6
XFILLER_0_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06075__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09800__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06075__B2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05822__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11206_ clknet_leaf_99_clk _00718_ net1166 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[678\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07575__A1 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11137_ clknet_leaf_86_clk _00649_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[609\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10841__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09316__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ clknet_leaf_41_clk _00580_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[540\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07327__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08524__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ net594 _01861_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_69_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10331__A0 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06535__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05889__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05984__S1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05560_ core.decoder.inst\[27\] _01392_ _01394_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08854__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10095__C1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05491_ _01588_ _01590_ net1030 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_60_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07230_ net989 core.register_file.registers_state\[577\] net875 core.register_file.registers_state\[609\]
+ net824 vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07161_ core.register_file.registers_state\[35\] core.register_file.registers_state\[3\]
+ net857 vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06066__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06112_ net939 core.register_file.registers_state\[808\] net759 net926 vssd1 vssd1
+ vccd1 vccd1 _02217_ sky130_fd_sc_hd__o31a_1
XANTENNA__07757__X _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07092_ _03195_ _03196_ net971 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11497__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06043_ net1037 core.register_file.registers_state\[138\] net668 core.register_file.registers_state\[170\]
+ net652 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07917__B _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07409__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05718__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout205 _04892_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08763__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout216 _04810_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
X_09802_ net560 _04834_ net459 net272 net1704 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__a32o_1
Xfanout238 net240 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
Xfanout249 _04690_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
X_07994_ _03748_ _03753_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__nand2_1
XANTENNA__06774__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _04938_ net297 net277 net2066 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__a22o_1
X_06945_ net987 core.register_file.registers_state\[715\] net864 core.register_file.registers_state\[747\]
+ net804 vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout280_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10322__A0 _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07869__A2 _03972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ net1107 core.register_file.registers_state\[142\] net847 core.register_file.registers_state\[174\]
+ net824 vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__o221a_1
X_09664_ _04806_ net295 net285 net2125 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__a22o_1
X_08615_ _04028_ _04243_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__or4_1
X_05827_ net940 core.register_file.registers_state\[656\] core.register_file.registers_state\[688\]
+ net697 net639 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a221o_1
X_09595_ _04955_ net403 net301 net2091 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout545_A _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1287_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ _04622_ _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__nand2_1
XANTENNA__08818__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05758_ net555 _01828_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09212__X _05031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08477_ core.pc.current_pc\[22\] net596 _04561_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_65_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08294__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05689_ net962 _01784_ _01785_ _01793_ net928 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a311oi_1
XANTENNA_fanout712_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06555__Y _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_X net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07428_ _03531_ _03532_ net1083 vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10714__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07359_ net1094 core.register_file.registers_state\[986\] core.register_file.registers_state\[1018\]
+ net835 net1071 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__o221a_1
XANTENNA__08046__A2 _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09243__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_X net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09794__A2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ net1539 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ net2005 net429 _04992_ net1002 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__a22o_1
XANTENNA__08930__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10864__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 net143 vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10253__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 core.register_file.registers_state\[302\] vssd1 vssd1 vccd1 vccd1 net1600
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 core.IO_mod.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05568__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout750 net752 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08939__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09534__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07843__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__buf_4
Xfanout772 _01468_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_107_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout783 _01462_ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_4
Xfanout794 _01455_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11237__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10313__A0 _05098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05363__A core.decoder.inst\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07190__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11824_ clknet_leaf_50_clk _01325_ net1307 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__dfrtp_1
XANTENNA__05740__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11755_ clknet_leaf_31_clk _00000_ net1206 vssd1 vssd1 vccd1 vccd1 core.ru.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06296__A1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10706_ clknet_leaf_69_clk _00218_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[178\]
+ sky130_fd_sc_hd__dfrtp_1
X_11686_ clknet_leaf_30_clk _01198_ net1201 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10637_ clknet_leaf_0_clk _00149_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09001__C _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload107 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06048__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07577__X _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09709__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09785__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10568_ clknet_leaf_95_clk _00080_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07796__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10499_ clknet_leaf_47_clk _00011_ net1291 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10163__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06220__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__X _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_1
X_06730_ net977 _02833_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__or3_1
XANTENNA__06369__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09170__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06661_ net1109 core.register_file.registers_state\[180\] net859 core.register_file.registers_state\[148\]
+ net814 vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07181__C1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ _02900_ _04335_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__o21ai_1
X_05612_ net939 core.register_file.registers_state\[695\] net749 net1011 vssd1 vssd1
+ vccd1 vccd1 _01717_ sky130_fd_sc_hd__o211a_1
X_09380_ net1768 net329 net321 _04791_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__a22o_1
X_06592_ net825 _02695_ _02696_ net786 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__o211a_1
XANTENNA__08584__A _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05560__X _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08331_ core.pc.current_pc\[9\] _04413_ core.pc.current_pc\[10\] vssd1 vssd1 vccd1
+ vccd1 _04428_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05543_ core.register_file.registers_state\[538\] net696 net638 _01647_ vssd1 vssd1
+ vccd1 vccd1 _01648_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_47_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08262_ core.pc.current_pc\[4\] _03260_ net577 vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05474_ net1043 core.register_file.registers_state\[477\] core.register_file.registers_state\[509\]
+ net672 net1011 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07213_ _03312_ _03317_ net781 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08193_ net530 _04288_ _04289_ _04297_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a31o_2
XANTENNA__08590__Y _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06039__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07144_ core.register_file.registers_state\[676\] core.register_file.registers_state\[644\]
+ net854 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10887__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__A _01987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09776__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08984__A0 _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07075_ core.register_file.registers_state\[742\] core.register_file.registers_state\[710\]
+ net839 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06026_ core.register_file.registers_state\[11\] net693 net636 _02130_ vssd1 vssd1
+ vccd1 vccd1 _02131_ sky130_fd_sc_hd__o211a_1
XANTENNA__05448__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10073__B net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07934__Y _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1202_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07977_ _03745_ _03777_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _04904_ net296 net276 net2525 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__a22o_1
X_06928_ net986 core.register_file.registers_state\[203\] net862 core.register_file.registers_state\[235\]
+ net802 vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09161__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _04707_ net296 net284 net2132 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__a22o_1
X_06859_ net538 _02052_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07172__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_36_clk_X clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ _04921_ net395 net299 net1695 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ _04607_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11540_ clknet_leaf_51_clk _01052_ net1297 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1012\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ clknet_leaf_83_clk _00983_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[943\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_135_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08941__B net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ net1407 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09767__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07778__A1 _03697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__C net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10353_ _05105_ net1549 net232 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05358__A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06450__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09519__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ net6 net902 net795 core.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__o22a_1
XANTENNA_input56_A gpio_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07844__Y _03949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09264__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout580 _03617_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
Xfanout591 net592 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_2
XFILLER_0_73_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11192__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07163__C1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11807_ clknet_leaf_52_clk _01308_ net1303 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09012__B _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11738_ clknet_leaf_47_clk _01250_ net1292 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08691__X _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06128__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09207__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ clknet_leaf_46_clk _01181_ net1291 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09758__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07900_ _03027_ _03402_ _03404_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_97_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08880_ net210 net2339 net372 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06729__C1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09391__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07831_ _03688_ _03927_ _03929_ _03931_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07762_ net531 _03866_ _03865_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_79_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09501_ net571 _04707_ net401 net309 net1657 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_49_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06713_ net1108 core.register_file.registers_state\[82\] core.register_file.registers_state\[114\]
+ net858 net813 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__o221a_1
X_07693_ net532 _03657_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__nand2_4
XFILLER_0_91_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06644_ _01827_ _02748_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__xnor2_1
X_09432_ net207 net738 net324 net313 net2137 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06827__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09363_ net1116 net463 _05021_ net413 net1672 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__a32o_1
X_06575_ core.register_file.registers_state\[279\] core.register_file.registers_state\[311\]
+ core.register_file.registers_state\[407\] core.register_file.registers_state\[439\]
+ net866 net1070 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout243_A _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ core.pc.current_pc\[8\] _04403_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__and2_1
X_05526_ net581 _01630_ _01628_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_30_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09294_ _04901_ net419 net333 net2324 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__a22o_1
XANTENNA__05468__C1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08245_ _04345_ _04348_ _04344_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_7_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05457_ core.register_file.registers_state\[541\] net696 net638 _01553_ vssd1 vssd1
+ vccd1 vccd1 _01562_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08761__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05877__S net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07658__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08176_ _01864_ net551 _03618_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09749__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05388_ _01408_ _01410_ core.decoder.inst\[31\] _01397_ vssd1 vssd1 vccd1 vccd1 _01493_
+ sky130_fd_sc_hd__and4b_1
XANTENNA__11065__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ _01632_ _02521_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08421__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06968__C1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1038_X net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07058_ net992 core.register_file.registers_state\[839\] net879 core.register_file.registers_state\[871\]
+ net1076 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a221o_1
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout877_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06009_ _02085_ _02113_ net582 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput194 net194 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XANTENNA__09382__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06291__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ clknet_leaf_19_clk _00483_ net1191 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[443\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08936__B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10259__A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_16_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07999__A1 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07999__B2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11408__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06175__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ clknet_leaf_65_clk _01035_ net1245 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[995\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06120__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05787__S _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06671__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11454_ clknet_leaf_94_clk _00966_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[926\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10405_ net1330 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11385_ clknet_leaf_60_clk _00897_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[857\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10336_ _05121_ net1606 net236 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__mux2_1
XANTENNA__05631__C1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__and2_1
XANTENNA__09373__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ net1126 net1498 net911 _05207_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__a31o_1
XANTENNA__07384__C1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07923__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05934__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09125__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08846__B _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10286__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05698__C1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09428__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10038__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06360_ net952 core.register_file.registers_state\[322\] net710 core.register_file.registers_state\[354\]
+ net1021 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_29_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05311_ core.control_logic.instruction\[6\] _01399_ net895 vssd1 vssd1 vccd1 vccd1
+ _01425_ sky130_fd_sc_hd__or3_1
XANTENNA__07749__Y _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06291_ core.register_file.registers_state\[291\] core.register_file.registers_state\[259\]
+ core.register_file.registers_state\[419\] core.register_file.registers_state\[387\]
+ net688 net1020 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06111__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08030_ _04025_ _04130_ _04134_ _03688_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput41 gpio_in[15] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput52 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold803 core.register_file.registers_state\[129\] vssd1 vssd1 vccd1 vccd1 net2122
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold814 core.register_file.registers_state\[617\] vssd1 vssd1 vccd1 vccd1 net2133
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 core.register_file.registers_state\[749\] vssd1 vssd1 vccd1 vccd1 net2144
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold836 core.register_file.registers_state\[377\] vssd1 vssd1 vccd1 vccd1 net2155
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold847 core.register_file.registers_state\[663\] vssd1 vssd1 vccd1 vccd1 net2166
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold858 core.register_file.registers_state\[834\] vssd1 vssd1 vccd1 vccd1 net2177
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09981_ _01421_ _01427_ net1315 vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold869 core.register_file.registers_state\[456\] vssd1 vssd1 vccd1 vccd1 net2188
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05622__C1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ net219 net739 vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05726__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _04795_ net2413 net374 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__mux2_1
XANTENNA__07914__B2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ _03538_ _03812_ _03512_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a21o_1
X_08794_ net606 net212 vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__and2_1
X_07745_ _01583_ _02630_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout360_A net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A _05060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08248__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06557__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ _03776_ _03780_ net484 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__mux2_1
XANTENNA__05689__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ net2327 net218 net406 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__mux2_1
XANTENNA__09419__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06627_ net783 _02723_ _02726_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__or3_1
XANTENNA__10079__A _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ net1119 _04990_ net414 net1612 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__a22o_1
X_06558_ net1094 core.register_file.registers_state\[983\] core.register_file.registers_state\[1015\]
+ net835 net1071 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__o221a_1
X_05509_ _01388_ _01403_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ net2524 net217 net338 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
X_06489_ net1035 core.register_file.registers_state\[472\] core.register_file.registers_state\[504\]
+ net670 net1009 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06653__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08228_ _03739_ _04332_ _04331_ _04328_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_132_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07850__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout994_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08159_ _01365_ _02052_ _02994_ _04263_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06405__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07602__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ clknet_leaf_78_clk _00682_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10121_ _05172_ _05173_ net588 vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09355__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ core.pc.current_pc\[1\] net589 vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__or2_1
XANTENNA__06231__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__C net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__C1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07118__C1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08666__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07570__B _03536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ clknet_leaf_106_clk _00466_ net1139 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[426\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07684__A3 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10885_ clknet_leaf_87_clk _00397_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09778__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09497__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11506_ clknet_leaf_65_clk _01018_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[978\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11437_ clknet_leaf_1_clk _00949_ net1139 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[909\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09594__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output87_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ clknet_leaf_13_clk _00880_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07745__B _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10319_ _05104_ net1817 net238 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08149__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ clknet_leaf_66_clk _00811_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[771\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09346__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05546__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09018__A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09897__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 net1153 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_2
Xfanout1161 net1167 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_4
X_05860_ net618 _01963_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__or3_1
XANTENNA__05907__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1172 net1179 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_2
Xfanout1183 net1184 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1196 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05791_ net1067 net897 _01867_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a21o_2
XANTENNA__07109__C1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07530_ _03633_ _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05281__A _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07461_ net632 _03565_ _03558_ net720 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a211o_2
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05712__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06332__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06412_ net586 _02514_ _02515_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09200_ _05005_ net358 net425 net1673 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__a22o_1
XANTENNA__05279__A_N core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07392_ core.register_file.registers_state\[537\] core.register_file.registers_state\[569\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06343_ net956 core.register_file.registers_state\[448\] net715 core.register_file.registers_state\[480\]
+ net930 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a221o_1
X_09131_ _04820_ net2518 net350 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08624__A2 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06383__Y _02488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09062_ net565 net603 net204 vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__and3_1
X_06274_ net634 _02378_ _01511_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11174__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08013_ net480 _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 core.register_file.registers_state\[616\] vssd1 vssd1 vccd1 vccd1 net1919
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout206_A _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold611 core.register_file.registers_state\[532\] vssd1 vssd1 vccd1 vccd1 net1930
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 core.register_file.registers_state\[614\] vssd1 vssd1 vccd1 vccd1 net1941
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold633 core.register_file.registers_state\[58\] vssd1 vssd1 vccd1 vccd1 net1952
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09585__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold644 core.register_file.registers_state\[264\] vssd1 vssd1 vccd1 vccd1 net1963
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06399__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold655 core.register_file.registers_state\[531\] vssd1 vssd1 vccd1 vccd1 net1974
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 core.register_file.registers_state\[387\] vssd1 vssd1 vccd1 vccd1 net1985
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 core.register_file.registers_state\[361\] vssd1 vssd1 vccd1 vccd1 net1996
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 core.register_file.registers_state\[225\] vssd1 vssd1 vccd1 vccd1 net2007
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07060__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ net1666 net2553 net798 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__mux2_1
XANTENNA__07655__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold699 core.register_file.registers_state\[85\] vssd1 vssd1 vccd1 vccd1 net2018
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1115_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ net567 _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__and2_1
XANTENNA__10081__B net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ net1115 _05073_ net378 net1629 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout575_A _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07348__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07899__B1 _04003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ _04655_ _04741_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__nor2_2
XANTENNA__08767__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05374__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ core.IO_mod.input_reg\[22\] net254 vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout742_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05989_ net1049 core.register_file.registers_state\[716\] vssd1 vssd1 vccd1 vccd1
+ _02094_ sky130_fd_sc_hd__or2_1
XANTENNA__05374__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07728_ _03639_ _03712_ net490 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__mux2_2
XANTENNA__07115__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ _03762_ _03763_ net484 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__mux2_2
XANTENNA__06323__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1272_X net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05677__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06874__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10670_ clknet_leaf_88_clk _00182_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[142\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08933__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09329_ net559 _04960_ _05052_ net332 net2472 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_11_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09576__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__B1_N _04179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09537__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ clknet_leaf_59_clk _00734_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[694\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08441__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07051__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07565__B _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ clknet_leaf_74_clk _00665_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[625\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05598__D1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09328__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ net1444 net516 _05161_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a21o_1
X_11084_ clknet_leaf_102_clk _00596_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[556\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ net724 _01611_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and2_2
XANTENNA__06896__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07581__A _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05460__S1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05532__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10937_ clknet_leaf_68_clk _00449_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[409\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08683__Y _04751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06865__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868_ clknet_leaf_51_clk _00380_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09803__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ clknet_leaf_83_clk _00311_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06078__C1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06617__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06617__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05825__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06712__S1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09567__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07042__A1 _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09319__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A2 _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06961_ _03062_ _03063_ _03065_ _03064_ net789 net816 vssd1 vssd1 vccd1 vccd1 _03066_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11276__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05707__C net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ net2038 net467 net434 _04765_ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__a22o_1
X_05912_ core.decoder.inst\[14\] net897 _01867_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__a21o_2
X_09680_ net207 net2301 net280 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06892_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08631_ core.decoder.inst\[7\] _04657_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05843_ _01946_ _01947_ net620 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ core.pc.current_pc\[30\] _04627_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__xnor2_1
X_05774_ _01877_ _01878_ net1028 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__o21a_1
XANTENNA__09098__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload95_A clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07513_ _01399_ _01499_ _01619_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__or3_4
X_08493_ _04556_ _04575_ _04565_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_18_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07444_ _02635_ _02662_ _03548_ _02633_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08526__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09211__A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__RESET_B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ _03478_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout323_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06608__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ _04730_ net2484 net350 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__mux2_1
XANTENNA__06608__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06326_ core.register_file.registers_state\[800\] core.register_file.registers_state\[768\]
+ core.register_file.registers_state\[928\] core.register_file.registers_state\[896\]
+ net692 net1022 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05816__C1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06257_ core.register_file.registers_state\[996\] core.register_file.registers_state\[964\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
X_09045_ _04659_ _04826_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__nor2_1
XANTENNA__07937__Y _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1232_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout209_X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06188_ net1044 core.register_file.registers_state\[486\] net750 _02292_ net924 vssd1
+ vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a311o_1
Xhold430 core.register_file.registers_state\[279\] vssd1 vssd1 vccd1 vccd1 net1749
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 core.register_file.registers_state\[785\] vssd1 vssd1 vccd1 vccd1 net1760
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 core.register_file.registers_state\[432\] vssd1 vssd1 vccd1 vccd1 net1771
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 core.register_file.registers_state\[267\] vssd1 vssd1 vccd1 vccd1 net1782
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold474 core.register_file.registers_state\[618\] vssd1 vssd1 vccd1 vccd1 net1793
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 core.CPU_DAT_I\[0\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1118_X net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold496 core.register_file.registers_state\[412\] vssd1 vssd1 vccd1 vccd1 net1815
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 _01449_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_4
Xfanout921 _01448_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_8
X_09947_ core.IO_mod.data_from_mem\[3\] core.CPU_DAT_O\[3\] net800 vssd1 vssd1 vccd1
+ vccd1 _01099_ sky130_fd_sc_hd__mux2_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_8
Xfanout943 _01374_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06792__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout954 net957 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06219__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout976 _01371_ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_8
Xfanout987 net997 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_4
X_09878_ _05053_ net459 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nand2_1
Xfanout998 _01368_ vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_8
Xhold1130 core.register_file.registers_state\[82\] vssd1 vssd1 vccd1 vccd1 net2449
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08533__A1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1141 core.register_file.registers_state\[600\] vssd1 vssd1 vccd1 vccd1 net2460
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05914__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09730__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08829_ net727 _03811_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__nand2_1
Xhold1152 core.register_file.registers_state\[116\] vssd1 vssd1 vccd1 vccd1 net2471
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1163 core.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_120_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 core.register_file.registers_state\[187\] vssd1 vssd1 vccd1 vccd1 net2493
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 core.register_file.registers_state\[458\] vssd1 vssd1 vccd1 vccd1 net2504
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 core.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ clknet_leaf_22_clk net66 net1181 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09820__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ clknet_leaf_24_clk _01275_ net1183 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10793__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__A2 _04878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__B net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10722_ clknet_leaf_77_clk _00234_ net1262 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[194\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10653_ clknet_leaf_17_clk _00165_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09797__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08960__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10584_ clknet_leaf_10_clk _00096_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload19 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_24_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07272__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09549__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09267__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05822__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10159__B2 core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11205_ clknet_leaf_100_clk _00717_ net1165 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07024__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08772__A1 _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11136_ clknet_leaf_58_clk _00648_ net1287 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[608\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11067_ clknet_leaf_21_clk _00579_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[539\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ net2305 net540 net519 _05109_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09015__B _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08827__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10095__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05490_ _01591_ _01592_ _01593_ _01594_ net622 net641 vssd1 vssd1 vccd1 vccd1 _01595_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08346__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09031__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07160_ net1111 core.register_file.registers_state\[131\] net857 core.register_file.registers_state\[163\]
+ net830 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__o221a_1
XANTENNA__09788__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10516__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06111_ net939 core.register_file.registers_state\[936\] net759 net1011 vssd1 vssd1
+ vccd1 vccd1 _02216_ sky130_fd_sc_hd__o31a_1
XANTENNA__07263__A1 _01372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07091_ net988 core.register_file.registers_state\[454\] net871 core.register_file.registers_state\[486\]
+ net980 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06042_ core.decoder.inst\[30\] net734 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__and2_1
XANTENNA__05558__X _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06471__C1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07015__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06449__S0 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10666__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout206 _04780_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06223__C1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout217 _04805_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09801_ net561 _04828_ net461 net272 net1780 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__a32o_1
Xfanout228 net231 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
X_07993_ _04078_ _04082_ net478 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload10_A clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ _04936_ net290 net275 net2362 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__a22o_1
X_06944_ net987 core.register_file.registers_state\[587\] net864 core.register_file.registers_state\[619\]
+ net816 vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09663_ _04801_ net286 net282 net2319 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06526__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ _02974_ _02977_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__o21a_1
X_08614_ _04064_ _04074_ _04268_ _04680_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__or4_1
XFILLER_0_136_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05826_ net1044 core.register_file.registers_state\[720\] core.register_file.registers_state\[752\]
+ net673 net654 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__o221a_1
X_09594_ _04953_ net396 net299 net2179 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08545_ _01551_ _04621_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nand2_1
X_05757_ _01853_ _01860_ net587 _01845_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_72_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08818__A2 _03964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ net231 _04556_ _04557_ _04560_ _04360_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__o32a_1
X_05688_ net948 core.register_file.registers_state\[1013\] net763 _01792_ net1029
+ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__o311a_1
XANTENNA__09491__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07427_ net1091 core.register_file.registers_state\[472\] core.register_file.registers_state\[504\]
+ net835 net1069 vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__o221a_1
XANTENNA__10087__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05501__A1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout705_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07358_ core.register_file.registers_state\[794\] core.register_file.registers_state\[826\]
+ core.register_file.registers_state\[922\] core.register_file.registers_state\[954\]
+ net866 net1071 vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux4_1
XANTENNA__08780__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07254__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06309_ net945 core.register_file.registers_state\[963\] vssd1 vssd1 vccd1 vccd1
+ _02414_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07289_ _03236_ _03393_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09794__A3 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1235_X net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ net745 net464 _04991_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07006__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 net166 vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 core.CPU_DAT_I\[16\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08779__X _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold282 core.register_file.registers_state\[269\] vssd1 vssd1 vccd1 vccd1 net1601
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07683__X _03788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10010__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 core.register_file.registers_state\[398\] vssd1 vssd1 vccd1 vccd1 net1612
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08939__B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 _04896_ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
Xfanout751 net752 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_2
Xfanout762 _01509_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_2
Xfanout773 _01468_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout784 net788 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09703__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout795 _05245_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_107_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06517__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07190__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09550__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11277__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ clknet_leaf_50_clk _01324_ net1308 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08809__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ clknet_leaf_30_clk net2114 net1202 vssd1 vssd1 vccd1 vccd1 wb.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06475__A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09482__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10705_ clknet_leaf_76_clk _00217_ net1260 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[177\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11528__SET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ clknet_leaf_31_clk _01197_ net1201 vssd1 vssd1 vccd1 vccd1 core.BUSY_O sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07858__X _03963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10636_ clknet_leaf_101_clk _00148_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09234__A2 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload108 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__inv_12
XANTENNA__07245__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10567_ clknet_leaf_92_clk _00079_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06453__C1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08993__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10498_ clknet_leaf_47_clk _00010_ net1306 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09942__A0 core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06205__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05559__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11119_ clknet_leaf_82_clk _00631_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[591\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05273__B core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06660_ net778 _02763_ _02764_ net774 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__o211a_1
XANTENNA__11314__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05611_ net1043 net749 core.register_file.registers_state\[663\] vssd1 vssd1 vccd1
+ vccd1 _01716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06591_ net993 core.register_file.registers_state\[662\] core.register_file.registers_state\[694\]
+ net880 net810 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a221o_1
XANTENNA__05731__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08330_ core.pc.current_pc\[9\] core.pc.current_pc\[10\] _04413_ vssd1 vssd1 vccd1
+ vccd1 _04427_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_47_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05542_ net939 core.register_file.registers_state\[570\] net759 vssd1 vssd1 vccd1
+ vccd1 _01647_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_47_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09473__A2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08261_ core.pc.current_pc\[3\] net598 _04364_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__o21ba_1
X_05473_ net1043 core.register_file.registers_state\[349\] core.register_file.registers_state\[381\]
+ net672 net925 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__o221a_1
XANTENNA__11464__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07484__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08681__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07212_ net1089 _03313_ _03316_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08192_ _03773_ _03866_ _04290_ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09225__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07143_ net778 _03241_ _03242_ net774 vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__B _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07074_ core.register_file.registers_state\[678\] core.register_file.registers_state\[646\]
+ net840 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__mux2_1
XANTENNA__05729__A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06025_ net936 core.register_file.registers_state\[43\] net760 vssd1 vssd1 vccd1
+ vccd1 _02130_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09528__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1028_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__A0 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A _05085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06211__A2 _02296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07976_ _03744_ _03747_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09715_ _04902_ net294 net276 net2143 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__a22o_1
X_06927_ net986 core.register_file.registers_state\[75\] net862 core.register_file.registers_state\[107\]
+ net816 vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout655_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09646_ _05022_ _05062_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__or2_4
X_06858_ _02084_ _02114_ _02526_ net538 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o31a_1
XFILLER_0_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07172__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05809_ _01911_ _01913_ net623 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a21o_1
X_09577_ _04919_ net395 net299 net1793 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06789_ net1097 core.register_file.registers_state\[592\] core.register_file.registers_state\[624\]
+ net839 net805 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ net593 _01665_ _04606_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__or3_1
XANTENNA__10269__A_N core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07475__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ _04543_ _04544_ _01782_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08427__B1_N net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ clknet_leaf_81_clk _00982_ net1235 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[942\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09216__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire448 _03629_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_1
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ net1339 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07227__B2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10352_ _05104_ net1585 net234 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__mux2_1
XANTENNA__06234__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07557__C _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08015__A _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06461__C net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ net5 net903 net795 core.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__o22a_1
XANTENNA__09924__A0 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09545__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input49_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06738__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06833__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11337__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 net573 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_4
Xfanout592 _05093_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08685__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09280__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11487__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06910__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11806_ clknet_leaf_54_clk _01307_ net1299 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09455__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07466__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11737_ clknet_leaf_46_clk _01249_ net1291 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__B2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11668_ clknet_leaf_46_clk _01180_ net1290 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06492__X _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09207__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10619_ clknet_leaf_23_clk _00131_ net1184 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11599_ clknet_leaf_24_clk _01111_ net1185 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08212__X _04317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08579__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ net489 _03934_ _03924_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ _03758_ _03770_ net491 vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__mux2_2
XANTENNA__05952__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05952__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ net1121 net605 _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__or3_4
XANTENNA__11128__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06712_ core.register_file.registers_state\[18\] core.register_file.registers_state\[50\]
+ core.register_file.registers_state\[146\] core.register_file.registers_state\[178\]
+ net889 net829 vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_49_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07692_ net510 _03658_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_49_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08595__A core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ _05026_ _05030_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__or2_4
X_06643_ _01865_ _02531_ net537 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05704__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05704__B2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09362_ net1117 net463 _05019_ net413 net1542 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__a32o_1
XANTENNA__10854__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06574_ net789 _02675_ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__o21a_1
XANTENNA__09446__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08313_ _04397_ _04401_ _04410_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a21oi_2
X_05525_ _01616_ _01620_ _01625_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__or3b_1
X_09293_ _04899_ net422 net333 net2046 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__a22o_1
XANTENNA__08654__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout236_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08244_ _04344_ _04345_ _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05456_ _01559_ _01560_ net959 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07209__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__C net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08175_ _01865_ _02779_ net548 net900 net1052 vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a32o_1
XANTENNA__05483__A3 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05387_ _01417_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout403_A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07126_ net769 _03217_ _03230_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__o21a_4
XFILLER_0_113_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07090__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07057_ net991 core.register_file.registers_state\[967\] net879 core.register_file.registers_state\[999\]
+ net983 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1312_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_105_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09906__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06008_ _02105_ _02112_ net722 _02097_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_A _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput195 net195 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1100_X net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07959_ net529 _04047_ _04062_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a21oi_4
XANTENNA__06291__S1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05943__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07556__A_N _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ clknet_leaf_9_clk _00482_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08936__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ net744 _05001_ net460 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09437__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08645__B1 _04716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05459__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07849__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07999__A2 _04100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ clknet_leaf_79_clk _01034_ net1253 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[994\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06120__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire245 _05246_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_134_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11453_ clknet_leaf_20_clk _00965_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[925\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_134_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ net1363 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11384_ clknet_leaf_3_clk _00896_ net1146 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[856\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10335_ _05120_ net1551 net238 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09275__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10266_ net2530 _05241_ _04360_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
XANTENNA__08399__B net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10727__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1310 net1311 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08176__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__S0 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ net68 net915 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__and2_1
XANTENNA__07384__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11221__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_X clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07136__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_41_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05310_ core.control_logic.instruction\[6\] net895 vssd1 vssd1 vccd1 vccd1 _01424_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06290_ net624 _02393_ _02394_ net634 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a31o_1
XFILLER_0_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06111__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_1
XFILLER_0_71_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput42 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput64 gpio_in[7] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
Xhold804 core.register_file.registers_state\[835\] vssd1 vssd1 vccd1 vccd1 net2123
+ sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_2
Xhold815 core.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 core.register_file.registers_state\[597\] vssd1 vssd1 vccd1 vccd1 net2145
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 core.register_file.registers_state\[495\] vssd1 vssd1 vccd1 vccd1 net2156
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold848 core.register_file.registers_state\[150\] vssd1 vssd1 vccd1 vccd1 net2167
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__A3 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ _01421_ _01427_ net1315 vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__o21ai_1
Xhold859 core.IO_mod.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ net2358 net369 _04927_ net436 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11652__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__RESET_B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ net220 net2283 net373 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__mux2_1
XANTENNA__08102__B _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _03512_ _03538_ _03812_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__nand3_1
XANTENNA__07914__A2 _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08793_ _04842_ _04843_ _04841_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__a21oi_4
XANTENNA__05925__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07470__S0 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07744_ net546 _03848_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09667__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05742__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__A1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout353_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ net2142 net219 net407 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
X_06626_ _02727_ _02728_ _02730_ _02729_ net786 net811 vssd1 vssd1 vccd1 vccd1 _02731_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10944__RESET_B net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06350__A1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10079__B net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06350__B2 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09345_ _04988_ net416 net412 net1652 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06557_ net553 _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout520_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_108_clk_X clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1262_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout618_A _01524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05508_ _01583_ _01612_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__or2_2
X_09276_ net2119 net218 net336 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
X_06488_ net1035 core.register_file.registers_state\[344\] core.register_file.registers_state\[376\]
+ net670 net923 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__o221a_1
XANTENNA__05536__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06573__A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08227_ _01499_ _01623_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07850__A1 _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05439_ net1047 core.register_file.registers_state\[350\] core.register_file.registers_state\[382\]
+ net674 net924 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05861__B1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ _02052_ _02994_ net578 vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout987_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ net989 core.register_file.registers_state\[709\] net875 core.register_file.registers_state\[741\]
+ net809 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__a221o_1
XANTENNA__07063__C1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ net487 _03721_ _03798_ _04189_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__o311a_1
X_10120_ net1124 core.pc.current_pc\[25\] core.pc.current_pc\[26\] vssd1 vssd1 vccd1
+ vccd1 _05173_ sky130_fd_sc_hd__or3_1
XANTENNA__07608__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08158__A2 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
X_10051_ net470 _05128_ _05129_ net516 net1498 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__a32o_1
XANTENNA__09823__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05916__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05377__C1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05916__B2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__B net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09658__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05652__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08866__A0 _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ clknet_leaf_16_clk _00465_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[425\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10884_ clknet_leaf_75_clk _00396_ net1262 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08963__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10614__RESET_B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09778__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05798__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07579__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06629__C1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ clknet_leaf_90_clk _01017_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[977\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11436_ clknet_leaf_103_clk _00948_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[908\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11367_ clknet_leaf_65_clk _00879_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[839\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ _05103_ net1560 net236 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__mux2_1
X_11298_ clknet_leaf_79_clk _00810_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[770\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09346__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ net86 net915 vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09018__B _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1140 net1179 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_2
Xfanout1151 net1153 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_4
Xfanout1162 net1167 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_2
XANTENNA__07452__S0 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05907__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1173 net1174 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_4
Xfanout1184 net1187 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
Xfanout1195 net1196 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_4
X_05790_ net582 _01893_ _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07109__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09649__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06580__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09034__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05281__B _01395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06868__C1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ _03560_ _03561_ _03563_ _03564_ net622 net645 vssd1 vssd1 vccd1 vccd1 _03565_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06332__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06411_ net586 _02514_ _02515_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_27_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07391_ core.register_file.registers_state\[729\] core.register_file.registers_state\[761\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08592__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_09130_ net215 net2359 net348 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06342_ net956 core.register_file.registers_state\[320\] net714 core.register_file.registers_state\[352\]
+ net1023 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_77_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06096__B1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09061_ net1773 net427 _05013_ net432 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06273_ net964 _02376_ _02377_ _02373_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08012_ net502 _03703_ _03698_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__o21a_1
XANTENNA__05843__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload40_A clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 core.register_file.registers_state\[281\] vssd1 vssd1 vccd1 vccd1 net1920
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold612 core.register_file.registers_state\[740\] vssd1 vssd1 vccd1 vccd1 net1931
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold623 core.register_file.registers_state\[773\] vssd1 vssd1 vccd1 vccd1 net1942
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09585__A1 _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 core.register_file.registers_state\[513\] vssd1 vssd1 vccd1 vccd1 net1953
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold645 core.register_file.registers_state\[34\] vssd1 vssd1 vccd1 vccd1 net1964
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06399__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10195__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold656 core.register_file.registers_state\[849\] vssd1 vssd1 vccd1 vccd1 net1975
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold667 core.register_file.registers_state\[425\] vssd1 vssd1 vccd1 vccd1 net1986
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ net1575 core.CPU_DAT_O\[19\] net800 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__mux2_1
Xhold678 core.register_file.registers_state\[367\] vssd1 vssd1 vccd1 vccd1 net1997
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08113__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__C _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 core.register_file.registers_state\[521\] vssd1 vssd1 vccd1 vccd1 net2008
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ _04763_ net602 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1010_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ net1118 _05072_ net376 net1751 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1108_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ _04736_ net2443 net373 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__mux2_1
XANTENNA__05359__C1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout470_A _05127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08767__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ net728 _04306_ _04757_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a21oi_1
X_05988_ core.register_file.registers_state\[748\] net675 vssd1 vssd1 vccd1 vccd1
+ _02093_ sky130_fd_sc_hd__or2_1
XANTENNA__06571__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06571__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07727_ net265 _03826_ _03827_ _03829_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout735_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_X net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ net497 _03719_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__or2_2
XANTENNA__06323__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06609_ net1105 core.register_file.registers_state\[470\] core.register_file.registers_state\[502\]
+ net852 net1080 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ _03616_ _03691_ _03693_ _02345_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_24_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05531__C1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09328_ core.register_file.registers_state\[383\] net475 net545 vssd1 vssd1 vccd1
+ vccd1 _05052_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09259_ _04882_ _05030_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__nor2_8
XFILLER_0_106_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07686__X _03791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ clknet_leaf_94_clk _00733_ net1242 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[693\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10186__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11152_ clknet_leaf_105_clk _00664_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[624\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ _04004_ net556 net589 core.pc.current_pc\[21\] net471 vssd1 vssd1 vccd1 vccd1
+ _05161_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_129_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11083_ clknet_leaf_108_clk _00595_ net1140 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[555\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07339__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ net1545 _05096_ net522 _05117_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08000__A1 _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07073__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10936_ clknet_leaf_10_clk _00448_ net1149 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[408\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06314__A1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08693__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08601__D_N _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07801__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10867_ clknet_leaf_12_clk _00379_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08980__X _04960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ clknet_leaf_89_clk _00310_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07596__X _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06093__A3 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09567__A1 _04899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ clknet_leaf_23_clk _00931_ net1184 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10177__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09319__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08790__A2 _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06250__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ core.register_file.registers_state\[938\] core.register_file.registers_state\[906\]
+ net832 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_05911_ net587 _02015_ _01989_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a21oi_4
XANTENNA_wire536_A _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07425__S0 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06891_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08630_ _04702_ _04703_ _04662_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a21oi_4
X_05842_ net1037 core.register_file.registers_state\[208\] core.register_file.registers_state\[240\]
+ net668 net652 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06553__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07750__B1 _03852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05292__A core.decoder.inst\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08561_ _04623_ _04635_ _04636_ _04637_ net228 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__a311oi_1
X_05773_ net1046 core.register_file.registers_state\[467\] core.register_file.registers_state\[499\]
+ net676 net1014 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07512_ _01399_ _01499_ _01619_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__nor3_4
X_08492_ _01747_ _04552_ _04566_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06305__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10101__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07443_ _03449_ net256 _03545_ _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__o31ai_4
XTAP_TAPCELL_ROW_18_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10595__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11840__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07374_ _03475_ _03477_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09255__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09211__B net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ _04724_ net2414 net350 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
XANTENNA__07266__C1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06325_ net1033 _02428_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09044_ net2401 net430 _05002_ net1001 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__a22o_1
X_06256_ core.register_file.registers_state\[932\] core.register_file.registers_state\[900\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07018__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 core.register_file.registers_state\[289\] vssd1 vssd1 vccd1 vccd1 net1739
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06187_ net940 core.register_file.registers_state\[454\] vssd1 vssd1 vccd1 vccd1
+ _02292_ sky130_fd_sc_hd__and2_1
Xhold431 core.register_file.registers_state\[771\] vssd1 vssd1 vccd1 vccd1 net1750
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10168__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1225_A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 core.register_file.registers_state\[570\] vssd1 vssd1 vccd1 vccd1 net1761
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold453 core.register_file.registers_state\[549\] vssd1 vssd1 vccd1 vccd1 net1772
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 core.register_file.registers_state\[410\] vssd1 vssd1 vccd1 vccd1 net1783
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 core.register_file.registers_state\[802\] vssd1 vssd1 vccd1 vccd1 net1794
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _01201_ vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10092__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout685_A _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout911 _01449_ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__buf_2
Xhold497 core.register_file.registers_state\[444\] vssd1 vssd1 vccd1 vccd1 net1816
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net926 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_4
X_09946_ core.IO_mod.data_from_mem\[2\] core.CPU_DAT_O\[2\] net800 vssd1 vssd1 vccd1
+ vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06792__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout933 _01375_ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net947 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net957 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout966 _01373_ vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06219__S1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout977 _01371_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1120 core.register_file.registers_state\[733\] vssd1 vssd1 vccd1 vccd1 net2439
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ net560 _04960_ net461 net268 net1664 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__a32o_1
Xfanout988 net997 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_4
Xfanout999 _01368_ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
Xhold1131 core.register_file.registers_state\[89\] vssd1 vssd1 vccd1 vccd1 net2450
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 core.register_file.registers_state\[723\] vssd1 vssd1 vccd1 vccd1 net2461
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08828_ core.IO_mod.data_from_mem\[30\] core.IO_mod.input_reg\[30\] net250 vssd1
+ vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__mux2_1
Xhold1153 core.register_file.registers_state\[383\] vssd1 vssd1 vccd1 vccd1 net2472
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10312__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1164 core.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06544__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07741__B1 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06544__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 core.register_file.registers_state\[81\] vssd1 vssd1 vccd1 vccd1 net2494
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 core.register_file.registers_state\[657\] vssd1 vssd1 vccd1 vccd1 net2505
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ net732 _04317_ net526 _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1197 core.register_file.registers_state\[209\] vssd1 vssd1 vccd1 vccd1 net2516
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11770_ clknet_leaf_24_clk _01274_ net1183 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09494__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10721_ clknet_leaf_88_clk _00233_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10652_ clknet_leaf_39_clk _00164_ net1218 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09246__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10267__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ clknet_leaf_20_clk _00095_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08960__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09548__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05902__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06480__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11204_ clknet_leaf_80_clk _00716_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[676\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07575__A3 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ clknet_leaf_40_clk _00647_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[607\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07980__A0 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__A _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ clknet_leaf_9_clk _00578_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[538\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ net724 _01893_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__and2_4
XANTENNA__05383__Y _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06535__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09485__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10095__A1 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07496__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ clknet_leaf_91_clk _00431_ net1239 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[391\]
+ sky130_fd_sc_hd__dfrtp_1
X_11899_ net1316 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06394__S0 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09031__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09237__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09788__A1 _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06110_ net1038 net749 core.register_file.registers_state\[904\] vssd1 vssd1 vccd1
+ vccd1 _02215_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07090_ net988 core.register_file.registers_state\[326\] net869 core.register_file.registers_state\[358\]
+ net1073 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11243__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06041_ _02117_ _02145_ net583 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_2
XFILLER_0_129_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08212__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06449__S1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08869__Y _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 _04705_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
X_09800_ net561 _04822_ net460 net271 net1879 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout218 _04800_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_2
Xfanout229 net230 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
X_07992_ _03115_ _04044_ _03086_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08598__A _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06774__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06774__B2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06943_ net816 _03046_ _03047_ net970 vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__o211a_1
X_09731_ _04934_ net296 net276 net2300 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__a22o_1
XANTENNA__10717__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05982__C1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _04796_ net295 net285 net1854 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06874_ net976 _02971_ _02978_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a21o_1
XANTENNA__06526__A1 _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__X _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ net255 _03811_ _04685_ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__or4_1
XANTENNA__07007__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05825_ net1044 core.register_file.registers_state\[592\] core.register_file.registers_state\[624\]
+ net673 net639 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__o221a_1
X_09593_ _04951_ net396 net299 net1945 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05734__C1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08544_ _01551_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05756_ _01853_ _01860_ _01845_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09476__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ _04558_ _04559_ net596 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout433_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05687_ net1054 core.register_file.registers_state\[981\] vssd1 vssd1 vccd1 vccd1
+ _01792_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1175_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07426_ net1091 core.register_file.registers_state\[344\] core.register_file.registers_state\[376\]
+ net835 net978 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09228__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10087__B net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07239__C1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07357_ net779 _03459_ _03461_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08780__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06308_ core.register_file.registers_state\[803\] core.register_file.registers_state\[771\]
+ core.register_file.registers_state\[931\] core.register_file.registers_state\[899\]
+ net687 net1020 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07288_ _03390_ _03391_ _03234_ _03264_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09027_ net614 net219 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__and2_1
X_06239_ core.decoder.inst\[25\] net734 net554 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1130_X net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 core.register_file.registers_state\[830\] vssd1 vssd1 vccd1 vccd1 net1569
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 net180 vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 _01217_ vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 core.ADR_I\[13\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06214__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 core.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__B2 _05105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net731 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_2
Xfanout741 _04655_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_6
XANTENNA__08939__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ net1066 net2455 net891 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
Xfanout752 net756 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05973__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_2
Xfanout774 _01468_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_4
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout785 net788 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_4
Xfanout796 _05245_ vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_107_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06517__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08020__B _03139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09831__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07190__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ clknet_leaf_49_clk _01323_ net1311 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11116__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09467__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11753_ clknet_leaf_31_clk _01265_ net1200 vssd1 vssd1 vccd1 vccd1 core.ru.prev_busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10704_ clknet_leaf_104_clk _00216_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[176\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ clknet_leaf_32_clk _01196_ net1206 vssd1 vssd1 vccd1 vccd1 core.SEL_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09219__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11266__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10635_ clknet_leaf_110_clk _00147_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09278__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_24_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ clknet_leaf_100_clk _00078_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08993__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10497_ net1362 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10881__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05559__A2 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06756__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11118_ clknet_leaf_90_clk _00630_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[590\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11049_ clknet_leaf_16_clk _00561_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[521\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XFILLER_0_56_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09170__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05273__C core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05610_ net939 core.register_file.registers_state\[567\] net759 vssd1 vssd1 vccd1
+ vccd1 _01715_ sky130_fd_sc_hd__or3_1
XANTENNA__09458__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06590_ core.register_file.registers_state\[534\] core.register_file.registers_state\[566\]
+ net880 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__mux2_1
XANTENNA__05731__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05541_ _01642_ _01645_ net721 _01640_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a211o_2
XANTENNA__11609__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08260_ net230 _04358_ _04359_ _04360_ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__o32a_1
XANTENNA__08681__A1 core.IO_mod.input_reg\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05472_ core.register_file.registers_state\[285\] core.register_file.registers_state\[317\]
+ core.register_file.registers_state\[413\] core.register_file.registers_state\[445\]
+ net696 net1011 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08881__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07211_ _03314_ _03315_ net976 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__a21o_1
XANTENNA__06692__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ _03864_ _03980_ _04291_ _04293_ _04295_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10633__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07142_ net1088 _03243_ _03246_ net781 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10240__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06444__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07073_ core.register_file.registers_state\[614\] core.register_file.registers_state\[582\]
+ net839 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__X _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06024_ net1036 core.register_file.registers_state\[139\] net667 core.register_file.registers_state\[171\]
+ net651 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05448__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07975_ _04078_ _04079_ net484 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__mux2_1
XANTENNA__06211__A3 _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06926_ _03028_ _03030_ net784 vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__o21a_1
X_09714_ _04900_ net292 net277 net2261 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__a22o_1
XANTENNA__09697__A0 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06857_ net769 _02961_ _02950_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__o21a_4
X_09645_ net567 _05062_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nor2_2
XANTENNA__07172__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1292_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05808_ core.register_file.registers_state\[18\] net690 net662 _01912_ vssd1 vssd1
+ vccd1 vccd1 _01913_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09576_ _04917_ net398 net302 net2133 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__a22o_1
X_06788_ net1097 core.register_file.registers_state\[720\] core.register_file.registers_state\[752\]
+ net839 net819 vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__o221a_1
XANTENNA__09449__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08527_ net593 _01665_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11289__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05739_ _01829_ _01832_ _01833_ net1032 net1006 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1080_X net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A _01460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ core.pc.current_pc\[21\] net574 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06132__C1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07409_ core.register_file.registers_state\[728\] core.register_file.registers_state\[760\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08389_ core.pc.current_pc\[15\] _02962_ net577 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ net1352 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10351_ _05103_ net1589 net232 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09826__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10282_ net4 net903 net795 net2550 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__o22a_1
XANTENNA__10639__RESET_B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__B1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__A1 core.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08727__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05655__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06833__S1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 net562 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_4
Xfanout571 net573 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_4
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_4
XANTENNA__09688__A0 _04887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout593 _01507_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08966__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07163__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06597__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11805_ clknet_leaf_72_clk _01306_ net1269 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11736_ clknet_leaf_46_clk _01248_ net1290 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09860__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05477__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11080__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ clknet_leaf_46_clk _01179_ net1290 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09207__A3 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10618_ clknet_leaf_5_clk _00130_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_11598_ clknet_leaf_26_clk _01110_ net1203 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09612__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10222__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10549_ clknet_leaf_63_clk _00061_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09915__A1 core.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06729__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07926__B1 _01958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07256__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__B2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09037__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06160__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05937__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ net511 _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__nand2_1
XANTENNA__08876__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ _02814_ _02815_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__nand2_1
XANTENNA__07780__A _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07691_ net265 _03791_ _03793_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_49_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08595__B _04656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09430_ net2287 net241 net406 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06642_ _02733_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__nor2_4
XANTENNA__06396__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09361_ _05017_ net418 net412 net1731 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__a22o_1
X_06573_ net784 _02676_ _02677_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__or3_1
XANTENNA__08103__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ _04397_ _04401_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__and3_1
XANTENNA__07779__X _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05524_ _01399_ _01415_ _01491_ _01622_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__nor4_1
XFILLER_0_129_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09292_ net1121 net601 _05030_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__or3_4
XANTENNA__08654__B2 _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_X clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05468__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08243_ _03382_ net575 _04346_ _02424_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a211oi_1
XANTENNA__05468__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06665__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05455_ net933 _01555_ _01556_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout229_A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ _02785_ _02905_ _03412_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05386_ net1003 _01366_ net896 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07125_ net777 _03224_ _03229_ net773 vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06968__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1138_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07090__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ core.register_file.registers_state\[807\] core.register_file.registers_state\[775\]
+ core.register_file.registers_state\[935\] core.register_file.registers_state\[903\]
+ net848 net1079 vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_06007_ net627 _02111_ net720 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1305_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput196 net196 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__09382__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05928__C1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07958_ _03925_ _03983_ _04002_ _04013_ net479 net495 vssd1 vssd1 vccd1 vccd1 _04063_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05762__X _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06909_ net1098 core.register_file.registers_state\[76\] core.register_file.registers_state\[108\]
+ net841 net806 vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__o221a_1
X_07889_ net513 _03992_ _03990_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09628_ net998 _05000_ net457 net391 net1711 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__a32o_1
XANTENNA__10320__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ net211 net1892 net305 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09842__A0 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05459__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ clknet_leaf_102_clk _01033_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[993\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_4_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11452_ clknet_leaf_41_clk _00964_ net1281 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[924\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_134_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06408__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ net1326 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11383_ clknet_leaf_22_clk _00895_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[855\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09556__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input61_A gpio_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _05119_ net1770 net239 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__mux2_1
XANTENNA__07865__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05631__B2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10265_ _04349_ _05240_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1300 net1301 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__clkbuf_4
Xfanout1311 net1312 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09373__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__S1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ net125 net917 net907 net1481 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__a22o_1
XANTENNA__07384__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05934__A2 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06768__X _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06592__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout390 _05085_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_4
XANTENNA__09291__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09144__X _05027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05490__S0 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05698__A1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09833__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11719_ clknet_leaf_49_clk net1568 net1309 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08207__Y _04312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06008__X _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
XFILLER_0_126_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput43 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput54 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05279__B core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput65 gpio_in[8] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold805 core.register_file.registers_state\[679\] vssd1 vssd1 vccd1 vccd1 net2124
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09061__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold816 core.register_file.registers_state\[757\] vssd1 vssd1 vccd1 vccd1 net2135
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold827 core.register_file.registers_state\[838\] vssd1 vssd1 vccd1 vccd1 net2146
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 core.register_file.registers_state\[674\] vssd1 vssd1 vccd1 vccd1 net2157
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07611__A2 _03289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold849 core.register_file.registers_state\[342\] vssd1 vssd1 vccd1 vccd1 net2168
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ net570 net220 net739 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__and3_1
XANTENNA__05622__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ _04890_ core.register_file.registers_state\[77\] net371 vssd1 vssd1 vccd1
+ vccd1 _00117_ sky130_fd_sc_hd__mux2_1
X_07812_ net527 _03886_ _03915_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07914__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05386__B1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08792_ core.IO_mod.input_reg\[24\] net250 net725 vssd1 vssd1 vccd1 vccd1 _04843_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07470__S1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ _01583_ _02630_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__nand2_1
XANTENNA__11349__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05481__S0 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07674_ _03777_ _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__nand2_1
XANTENNA__07678__A2 _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05689__A1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ net2264 net220 net407 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
X_06625_ core.register_file.registers_state\[853\] core.register_file.registers_state\[885\]
+ net879 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XANTENNA__06886__B1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout346_A _05027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06556_ _01612_ _02601_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__xor2_1
XANTENNA__09824__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ net1115 net463 _04986_ net413 net1520 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05507_ _01585_ _01611_ net582 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07835__C1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09275_ net2240 net219 net337 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
X_06487_ net958 _02591_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout513_A _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10984__RESET_B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05536__S1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ _03738_ _04326_ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05438_ core.register_file.registers_state\[286\] core.register_file.registers_state\[318\]
+ core.register_file.registers_state\[414\] core.register_file.registers_state\[446\]
+ net703 net1017 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07850__A2 _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10913__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08157_ _02052_ _02994_ _03621_ _02017_ net900 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05369_ net1084 _01470_ _01473_ net780 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_X net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09052__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07108_ net989 core.register_file.registers_state\[581\] net875 core.register_file.registers_state\[613\]
+ net824 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a221o_1
XANTENNA__07602__A2 _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ _03622_ _04190_ _04191_ _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout882_A _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05613__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07039_ _03142_ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1210_X net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ _04242_ net588 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__nand2_1
XANTENNA__09355__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07366__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05472__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05933__A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10122__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10952_ clknet_leaf_12_clk _00464_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[424\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10883_ clknet_leaf_73_clk _00395_ net1272 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[355\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08963__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08079__C1 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__A0 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06629__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07579__B _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09291__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11504_ clknet_leaf_103_clk _01016_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[976\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_109_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05852__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11435_ clknet_leaf_108_clk _00947_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[907\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10189__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09286__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ clknet_leaf_105_clk _00878_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[838\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08043__X _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ _05102_ net1461 net236 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11297_ clknet_leaf_85_clk _00809_ net1236 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10844__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10248_ net1125 net1436 net911 _05232_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_33_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07357__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1130 net1134 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_4
Xfanout1141 net1142 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10361__A0 _05113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__clkbuf_4
X_10179_ net106 net917 net907 net2495 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__a22o_1
Xfanout1163 net1166 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06565__C1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07452__S1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1174 net1178 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07534__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1185 net1186 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_4
Xfanout1196 net1202 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_2
XFILLER_0_117_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07109__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09034__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06410_ net586 _02488_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07390_ core.register_file.registers_state\[665\] core.register_file.registers_state\[697\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
XANTENNA__06674__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05540__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06341_ net1032 _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09282__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09060_ net565 _05012_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06272_ net929 _02375_ net1031 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08011_ _04025_ _04037_ _04113_ net547 _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold602 core.register_file.registers_state\[470\] vssd1 vssd1 vccd1 vccd1 net1921
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold613 core.register_file.registers_state\[612\] vssd1 vssd1 vccd1 vccd1 net1932
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 core.register_file.registers_state\[516\] vssd1 vssd1 vccd1 vccd1 net1943
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09585__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold635 core.register_file.registers_state\[533\] vssd1 vssd1 vccd1 vccd1 net1954
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 core.register_file.registers_state\[613\] vssd1 vssd1 vccd1 vccd1 net1965
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold657 core.register_file.registers_state\[569\] vssd1 vssd1 vccd1 vccd1 net1976
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold668 core.register_file.registers_state\[554\] vssd1 vssd1 vccd1 vccd1 net1987
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net1618 core.CPU_DAT_O\[18\] net798 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__mux2_1
Xhold679 core.register_file.registers_state\[856\] vssd1 vssd1 vccd1 vccd1 net1998
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08888__X _04899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__D net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09337__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08913_ core.register_file.registers_state\[104\] net368 _04915_ net434 vssd1 vssd1
+ vccd1 vccd1 _00144_ sky130_fd_sc_hd__a22o_1
X_09893_ net1118 _05071_ net376 net1852 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07348__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__A0 _05104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ net224 net2478 net373 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1003_A _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08767__C net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05987_ net1049 core.register_file.registers_state\[588\] core.register_file.registers_state\[620\]
+ net675 net639 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__o221a_1
X_08775_ net2147 net468 net437 _04828_ vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout463_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11112__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ net498 _03659_ _03825_ _03830_ net490 vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07657_ _03760_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout630_A _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ net1105 core.register_file.registers_state\[342\] core.register_file.registers_state\[374\]
+ net851 net985 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__o221a_1
XANTENNA__08275__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07588_ net1114 _01407_ _01417_ _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06539_ net975 _02642_ _02643_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__or3_1
X_09327_ _04959_ net417 net332 net2016 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a22o_1
XANTENNA__10717__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1160_X net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09258_ net560 _04881_ _05045_ net340 net2094 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_131_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08209_ net1114 _04311_ _04313_ net580 vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_116_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07871__A1_N net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09189_ _04983_ net351 net423 net1782 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_116_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11220_ clknet_leaf_55_clk _00732_ net1295 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[692\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07619__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ clknet_leaf_79_clk _00663_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[623\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08798__X _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05598__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net1454 net516 _05160_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_129_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09834__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09328__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ clknet_leaf_106_clk _00594_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[554\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07339__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _01688_ _01706_ net724 vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_125_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10343__A0 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06011__A1 core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06011__B2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10935_ clknet_leaf_21_clk _00447_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[407\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07824__A1_N core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ clknet_leaf_68_clk _00378_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[338\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09264__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ clknet_leaf_2_clk _00309_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06078__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09803__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07275__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06078__B2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05825__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05825__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output92_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11792__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ clknet_leaf_6_clk _00930_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[890\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06433__S net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08214__A _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07578__A1 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08775__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11349_ clknet_leaf_62_clk _00861_ net1242 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06786__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05910_ net718 _02014_ _02003_ _01995_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA_clkbuf_leaf_107_clk_X clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06890_ _02052_ _02963_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06538__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07425__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05573__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05841_ net1037 core.register_file.registers_state\[80\] core.register_file.registers_state\[112\]
+ net668 net637 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09045__A _04659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08560_ _04623_ _04636_ _04635_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a21oi_1
X_05772_ net1050 core.register_file.registers_state\[339\] core.register_file.registers_state\[371\]
+ net676 net924 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__o221a_1
XANTENNA__05761__B1 _01862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07511_ _01366_ _01400_ _01429_ _01622_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__or4_4
XFILLER_0_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08491_ _02562_ _04572_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06936__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07442_ _02662_ _03546_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10576__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07373_ _03475_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06324_ net955 core.register_file.registers_state\[576\] net713 core.register_file.registers_state\[608\]
+ net662 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a221o_1
X_09112_ net226 net2314 net349 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07266__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06069__B2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08823__S net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05816__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09043_ net744 net464 _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06255_ core.register_file.registers_state\[868\] core.register_file.registers_state\[836\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout211_A _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold410 net111 vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06186_ net1044 core.register_file.registers_state\[358\] net750 _02290_ vssd1 vssd1
+ vccd1 vccd1 _02291_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold421 net187 vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 core.register_file.registers_state\[911\] vssd1 vssd1 vccd1 vccd1 net1751
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 core.register_file.registers_state\[423\] vssd1 vssd1 vccd1 vccd1 net1762
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold454 core.register_file.registers_state\[154\] vssd1 vssd1 vccd1 vccd1 net1773
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold465 core.register_file.registers_state\[703\] vssd1 vssd1 vccd1 vccd1 net1784
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A core.decoder.inst\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold476 core.register_file.registers_state\[159\] vssd1 vssd1 vccd1 vccd1 net1795
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06241__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1218_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 core.register_file.registers_state\[290\] vssd1 vssd1 vccd1 vccd1 net1806
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _01396_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_2
Xhold498 net176 vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout912 _01449_ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09945_ core.IO_mod.data_from_mem\[1\] core.CPU_DAT_O\[1\] net799 vssd1 vssd1 vccd1
+ vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout580_A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 net926 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout934 _01375_ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_6
XFILLER_0_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net946 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10325__A0 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_2
Xfanout967 _01372_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _04959_ net390 net268 net2159 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11515__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout978 net981 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__buf_4
Xhold1110 core.register_file.registers_state\[115\] vssd1 vssd1 vccd1 vccd1 net2429
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net990 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09191__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1121 core.register_file.registers_state\[371\] vssd1 vssd1 vccd1 vccd1 net2440
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 core.register_file.registers_state\[101\] vssd1 vssd1 vccd1 vccd1 net2451
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09730__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08827_ net2182 net466 net462 _04872_ vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__a22o_1
Xhold1143 core.register_file.registers_state\[577\] vssd1 vssd1 vccd1 vccd1 net2462
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05914__C net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 core.register_file.registers_state\[654\] vssd1 vssd1 vccd1 vccd1 net2473
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1165 core.register_file.registers_state\[195\] vssd1 vssd1 vccd1 vccd1 net2484
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_120_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1176 core.CPU_DAT_I\[14\] vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 core.register_file.registers_state\[97\] vssd1 vssd1 vccd1 vccd1 net2506
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ core.IO_mod.data_from_mem\[19\] net247 _04813_ vssd1 vssd1 vccd1 vccd1 _04814_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08794__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1198 core.register_file.registers_state\[136\] vssd1 vssd1 vccd1 vccd1 net2517
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_105_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _03543_ _03812_ _03480_ _03510_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__a211o_1
X_08689_ _04700_ _04718_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09494__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ clknet_leaf_52_clk _00232_ net1302 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[192\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06701__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06518__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08049__A2 _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ clknet_leaf_23_clk _00163_ net1186 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09829__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09797__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ clknet_leaf_59_clk _00094_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08960__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05902__S1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11045__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11203_ clknet_leaf_67_clk _00715_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[675\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ clknet_leaf_95_clk _00646_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[606\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05440__C1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__B _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10316__A0 _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11065_ clknet_leaf_68_clk _00577_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[537\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07084__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ net1485 net542 net521 _05108_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__a22o_1
XANTENNA__09182__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09721__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07193__C1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06091__S0 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05743__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10095__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ clknet_leaf_101_clk _00430_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[390\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11898_ net100 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06394__S1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09237__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10849_ clknet_leaf_86_clk _00361_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[321\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09788__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06040_ net717 _02128_ _02136_ _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__o22a_4
XANTENNA__06471__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06471__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11538__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06223__A1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout208 _04334_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08231__X _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout219 _04795_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
X_07991_ net528 _04076_ _04077_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o211a_2
XFILLER_0_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08598__B _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _04932_ net294 net276 net2107 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__a22o_1
X_06942_ net1093 core.register_file.registers_state\[683\] core.register_file.registers_state\[651\]
+ net833 net804 vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a221o_1
XANTENNA__10307__A0 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05507__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09661_ _04791_ net295 net284 net2076 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__a22o_1
X_06873_ net1088 _02969_ _02970_ net967 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08612_ _03839_ _04672_ _04686_ _03964_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__or4b_1
X_05824_ net585 _01927_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__or2_1
X_09592_ _04949_ net402 net301 net1910 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__a22o_1
XANTENNA__06931__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08543_ core.pc.current_pc\[29\] _02630_ net574 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__mux2_1
X_05755_ net630 _01859_ net718 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout259_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__X _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ core.pc.current_pc\[22\] _04540_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05686_ net1056 core.register_file.registers_state\[853\] vssd1 vssd1 vccd1 vccd1
+ _01791_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07425_ core.register_file.registers_state\[280\] core.register_file.registers_state\[312\]
+ core.register_file.registers_state\[408\] core.register_file.registers_state\[440\]
+ net865 net1072 vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07239__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ net969 _03452_ _03460_ net775 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06862__A _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08987__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06307_ net964 _02405_ _02406_ _02411_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a31o_1
X_07287_ _03390_ _03391_ _03264_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ net2489 net429 _04990_ net1002 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__a22o_1
X_06238_ _02335_ _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__and2_4
XANTENNA__06462__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08739__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06169_ core.decoder.inst\[27\] net734 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__nand2_1
Xhold240 net167 vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09400__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 core.register_file.registers_state\[46\] vssd1 vssd1 vccd1 vccd1 net1570
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold262 core.CPU_DAT_I\[6\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 core.register_file.registers_state\[528\] vssd1 vssd1 vccd1 vccd1 net1592
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10010__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 core.IO_mod.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 core.IO_mod.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout962_A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout720 _01512_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_6
XANTENNA__05568__A3 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07962__B2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 _01420_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10323__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09928_ net1071 core.CPU_DAT_O\[17\] net891 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
Xfanout742 net746 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
Xfanout753 net756 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_4
Xfanout764 net766 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07980__X _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09164__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout775 _01463_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout786 net787 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout797 _05244_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_2
XANTENNA__06102__A core.decoder.inst\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _04925_ net383 net266 net1819 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__a22o_1
XANTENNA__07175__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07632__S net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05941__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ clknet_leaf_47_clk _01322_ net1292 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11752_ clknet_leaf_31_clk _01264_ net1206 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06248__S net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10703_ clknet_leaf_84_clk _00215_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[175\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11683_ clknet_leaf_32_clk _01195_ net1205 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08971__B net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09559__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ clknet_leaf_111_clk _00146_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07325__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10565_ clknet_leaf_96_clk _00077_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07079__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06453__A1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11286__RESET_B net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10496_ net1401 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11215__RESET_B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08699__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05675__X _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07402__B1 _02534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05559__A3 _01663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05413__C1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ clknet_leaf_4_clk _00629_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[589\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09155__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ clknet_leaf_12_clk _00560_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[520\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
XFILLER_0_95_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06913__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wire227_A _04719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05540_ net958 _01643_ _01644_ net631 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__o31a_1
XFILLER_0_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07469__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06158__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08130__A1 _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05471_ _01572_ _01575_ _01521_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11210__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06141__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07210_ net994 core.register_file.registers_state\[450\] net884 core.register_file.registers_state\[482\]
+ net983 vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__a221o_1
X_08190_ net1112 _04292_ _04294_ net578 vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__o211a_1
XANTENNA__06692__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07141_ _03244_ _03245_ net976 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08433__A2 _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05298__A core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07072_ core.register_file.registers_state\[550\] core.register_file.registers_state\[518\]
+ net840 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__mux2_1
XANTENNA__05878__S0 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05729__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06023_ _02122_ _02127_ net631 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XANTENNA__10928__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08197__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09394__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07974_ net506 _03632_ _03785_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a21o_1
XANTENNA__05955__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09713_ net207 net738 net296 net276 net1864 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__a32o_1
X_06925_ core.register_file.registers_state\[11\] net864 net802 _03029_ vssd1 vssd1
+ vccd1 vccd1 _03030_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout376_A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ net999 _05021_ net457 net392 net1737 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__a32o_1
X_06856_ _02955_ _02960_ net781 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__mux2_1
X_05807_ net1060 core.register_file.registers_state\[50\] net755 vssd1 vssd1 vccd1
+ vccd1 _01912_ sky130_fd_sc_hd__and3_1
X_09575_ _04915_ net397 net302 net1919 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout543_A _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06787_ net971 _02890_ _02891_ net1067 vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout1285_A net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08526_ core.pc.current_pc\[27\] _03446_ net574 vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05738_ _01835_ _01838_ _01839_ _01842_ net934 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_19_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08457_ _02747_ net575 vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__nand2_1
XANTENNA__07959__Y _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05669_ net949 core.register_file.registers_state\[502\] net764 _01773_ net1022 vssd1
+ vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07408_ core.register_file.registers_state\[664\] core.register_file.registers_state\[696\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07880__B1 _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ core.pc.current_pc\[15\] _04477_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07339_ net969 _03442_ _03443_ net1066 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__o31a_1
XANTENNA__10318__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09621__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _05102_ net1492 net232 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09009_ net604 _04888_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__and2_1
XANTENNA__11853__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10281_ net3 net904 net797 core.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__B2 _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09385__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06738__A2 _01987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09842__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout572 net573 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_4
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_2
XANTENNA__10608__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 _01502_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_8
XANTENNA__07870__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06597__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11804_ clknet_leaf_52_clk _01305_ net1303 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08982__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11735_ clknet_leaf_46_clk _01247_ net1289 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09289__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ clknet_leaf_46_clk _01178_ net1289 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07871__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10617_ clknet_leaf_70_clk _00129_ net1275 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_11597_ clknet_leaf_29_clk _01109_ net1200 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08206__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10548_ clknet_leaf_54_clk _00060_ net1300 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10479_ net1487 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08179__A1 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__B2 _03950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09376__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05846__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06441__S net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A1 _01987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__B2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09037__B net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05937__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09128__A0 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07139__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08876__B _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ net550 _02813_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07780__B _03422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ net1112 _03792_ _03794_ net580 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__o211a_1
XANTENNA__06677__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09053__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ net783 _02744_ _02745_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09360_ net1116 _05016_ net413 net1815 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10600__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06572_ net1095 core.register_file.registers_state\[215\] core.register_file.registers_state\[247\]
+ net836 net818 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__o221a_1
XANTENNA__08103__A1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08311_ _04408_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__or2_1
XANTENNA__09300__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05523_ _01615_ _01626_ _01627_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__o21a_1
X_09291_ net2419 net241 net336 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
XANTENNA__08654__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08242_ _03382_ net575 vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__and2_1
X_05454_ net1005 _01557_ _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__or3_1
XANTENNA__09500__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05295__C_N core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05873__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ _04270_ _04271_ _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__and3_4
X_05385_ _01417_ _01489_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__or2_2
XANTENNA__11876__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09603__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09927__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ net1086 _03225_ _03228_ net783 vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07090__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ _03151_ _03154_ _03159_ net769 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o211a_1
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
X_06006_ net1027 _02109_ _02110_ _02106_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__o22a_1
XANTENNA__09367__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XANTENNA__09906__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__07378__C1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
Xoutput197 net197 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10772__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__A0 _04887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06196__A3 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07957_ net265 _04060_ _04061_ _04048_ _04053_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__a2111o_2
XANTENNA_fanout660_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ net1098 core.register_file.registers_state\[204\] core.register_file.registers_state\[236\]
+ net841 net820 vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07888_ net513 _03992_ _03990_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ net2497 net393 _05075_ net1001 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06839_ net1107 core.register_file.registers_state\[143\] net847 core.register_file.registers_state\[175\]
+ net826 vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1190_X net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09558_ net212 net2460 net303 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08509_ _04590_ _04584_ net228 vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08645__A2 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ _05008_ net317 net261 net1856 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ clknet_leaf_58_clk _01032_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[992\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07853__B1 _03956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11560__RESET_B net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05864__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11451_ clknet_leaf_22_clk _00963_ net1181 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[923\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06408__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ net1346 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09837__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11382_ clknet_leaf_42_clk _00894_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[854\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05616__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10333_ _05118_ net1753 net239 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05666__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09358__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ _04344_ _04345_ _04348_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__a21oi_1
Xfanout1301 net1305 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__buf_2
X_10195_ net124 net919 net909 net1567 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__a22o_1
Xfanout1312 net1313 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__buf_2
XANTENNA__08977__A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05490__S1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08333__A1 _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06344__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11718_ clknet_leaf_49_clk net1596 net1310 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06436__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06111__A3 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11649_ clknet_leaf_49_clk _01161_ net1310 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09597__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_1
Xinput44 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput55 gpio_in[28] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09061__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput66 gpio_in[9] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold806 core.register_file.registers_state\[689\] vssd1 vssd1 vccd1 vccd1 net2125
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold817 core.register_file.registers_state\[903\] vssd1 vssd1 vccd1 vccd1 net2136
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold828 core.register_file.registers_state\[53\] vssd1 vssd1 vccd1 vccd1 net2147
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 core.register_file.registers_state\[610\] vssd1 vssd1 vccd1 vccd1 net2158
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09349__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09048__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11279__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06258__S0 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08860_ net741 _04785_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nor2_2
XANTENNA__08887__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ net527 _03886_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__o21a_1
XANTENNA__05386__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08791_ core.IO_mod.data_from_mem\[24\] net246 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__nand2_1
X_07742_ _03665_ _03673_ _03845_ net493 _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__o221a_1
XANTENNA__05481__S1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__A1 core.decoder.inst\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09521__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ net452 _02900_ net444 net501 vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a31o_1
XANTENNA__06335__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05742__C net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__A3 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09412_ net2404 _04890_ net405 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06624_ core.register_file.registers_state\[789\] core.register_file.registers_state\[821\]
+ net879 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09343_ net1115 _04984_ net412 net2196 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__a22o_1
X_06555_ net553 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__inv_2
XANTENNA__08627__A2 _03739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_A _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_A _05031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05506_ net723 _01598_ _01603_ _01610_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__o22a_1
X_09274_ net2175 net220 net337 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08127__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06486_ core.register_file.registers_state\[280\] core.register_file.registers_state\[312\]
+ core.register_file.registers_state\[408\] core.register_file.registers_state\[440\]
+ net695 net1009 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08225_ _04324_ _04327_ _04329_ net255 vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05437_ _01538_ _01541_ net632 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1150_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1248_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ _02935_ _02998_ _04005_ net530 vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__o31a_1
X_05368_ net971 _01471_ _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__or3_1
XANTENNA__10198__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09052__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ net819 _03210_ _03211_ net974 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__o211a_1
XANTENNA__07063__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08260__B1 _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05757__Y _01862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05299_ core.decoder.inst\[27\] core.decoder.inst\[28\] core.decoder.inst\[29\] vssd1
+ vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__or3_1
X_08087_ net533 _03290_ _03618_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07177__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07038_ _03111_ _03114_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__nand2_1
XANTENNA__06081__S net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__B2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08563__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09760__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05377__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net743 net465 _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05377__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05472__S1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09512__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ clknet_leaf_92_clk _00463_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[423\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05652__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10122__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10882_ clknet_leaf_78_clk _00394_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[354\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08963__C net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11059__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06629__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06256__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ clknet_leaf_79_clk _01015_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[975\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09579__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07876__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05852__A2 _01956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ clknet_leaf_107_clk _00946_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[906\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06780__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07054__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11365_ clknet_leaf_86_clk _00877_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[837\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_100_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05396__A _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10316_ _05101_ net1978 net238 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11296_ clknet_leaf_56_clk _00808_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[768\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10247_ net85 net914 vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1120 core.decoder.inst\[10\] vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_4
Xfanout1131 net1134 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09751__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1142 net1146 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1153 net1179 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_2
X_10178_ net105 net917 net907 net1587 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__a22o_1
Xfanout1164 net1166 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1175 net1177 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_4
Xfanout1186 net1187 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_2
Xfanout1197 net1202 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08306__B2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09503__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06868__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06868__B2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05540__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06340_ core.register_file.registers_state\[288\] core.register_file.registers_state\[256\]
+ core.register_file.registers_state\[416\] core.register_file.registers_state\[384\]
+ net691 net1022 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06271_ core.register_file.registers_state\[292\] core.register_file.registers_state\[260\]
+ core.register_file.registers_state\[420\] core.register_file.registers_state\[388\]
+ net688 net1021 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08010_ net1113 _04113_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold603 core.register_file.registers_state\[906\] vssd1 vssd1 vccd1 vccd1 net1922
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold614 core.register_file.registers_state\[507\] vssd1 vssd1 vccd1 vccd1 net1933
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold625 core.register_file.registers_state\[758\] vssd1 vssd1 vccd1 vccd1 net1944
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold636 core.register_file.registers_state\[750\] vssd1 vssd1 vccd1 vccd1 net1955
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold647 core.register_file.registers_state\[362\] vssd1 vssd1 vccd1 vccd1 net1966
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold658 core.ADR_I\[29\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06253__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09961_ net1583 core.CPU_DAT_O\[17\] net798 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__mux2_1
XANTENNA__09990__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold669 core.register_file.registers_state\[813\] vssd1 vssd1 vccd1 vccd1 net1988
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload26_A clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ net567 _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09892_ _04988_ net383 net375 net1855 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__a22o_1
XANTENNA__09742__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _04724_ net2447 net373 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__mux2_1
XANTENNA__05359__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05359__B2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout289_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ net570 _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05986_ net941 core.register_file.registers_state\[652\] core.register_file.registers_state\[684\]
+ net698 net640 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a221o_1
XANTENNA__09940__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07725_ _03821_ _03822_ net483 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06859__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06403__S0 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ net500 net449 _03320_ net441 vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06607_ core.register_file.registers_state\[278\] core.register_file.registers_state\[310\]
+ core.register_file.registers_state\[406\] core.register_file.registers_state\[438\]
+ net880 net1080 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05531__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _01400_ _01493_ _01617_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout623_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05531__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09326_ _04957_ net418 net332 net2050 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06538_ net1104 core.register_file.registers_state\[476\] core.register_file.registers_state\[508\]
+ net852 net1077 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09257_ core.register_file.registers_state\[319\] net475 _04708_ vssd1 vssd1 vccd1
+ vccd1 _05045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06469_ net1004 _02570_ _02573_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08208_ _01895_ net550 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ _04981_ net351 net423 net1640 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__a22o_1
XANTENNA__06804__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08139_ _03957_ _04089_ net531 vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10040__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11150_ clknet_leaf_90_clk _00662_ net1235 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[622\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _04287_ net557 net589 core.pc.current_pc\[20\] net471 vssd1 vssd1 vccd1 vccd1
+ _05160_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_129_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11081_ clknet_leaf_16_clk _00593_ net1216 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[553\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09733__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ net2481 net541 net520 _05116_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05770__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08974__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10934_ clknet_leaf_60_clk _00446_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[406\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08466__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06775__A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ clknet_leaf_72_clk _00377_ net1272 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10796_ clknet_leaf_102_clk _00308_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10811__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06483__C1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07027__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05397__Y _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11417_ clknet_leaf_56_clk _00929_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08214__B _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ clknet_leaf_56_clk _00860_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[820\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05589__A1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06250__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ clknet_leaf_82_clk _00791_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[751\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07545__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08527__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09724__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05840_ net652 _01944_ _01943_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09045__B _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A2 _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05771_ core.register_file.registers_state\[275\] core.register_file.registers_state\[307\]
+ core.register_file.registers_state\[403\] core.register_file.registers_state\[435\]
+ net697 net1014 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05761__A1 _01825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07510_ _02604_ _03550_ _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07189__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08490_ _02562_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__and2b_1
XANTENNA__08376__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06305__A3 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06936__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07441_ net553 _02661_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07372_ _01664_ _02600_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09255__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ _04704_ net2454 net349 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07266__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06323_ net955 core.register_file.registers_state\[704\] net713 core.register_file.registers_state\[736\]
+ net648 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09042_ net613 net214 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__and2_1
X_06254_ core.register_file.registers_state\[804\] core.register_file.registers_state\[772\]
+ net687 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06624__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07018__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold400 core.register_file.registers_state\[305\] vssd1 vssd1 vccd1 vccd1 net1719
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07018__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06185_ net940 core.register_file.registers_state\[326\] net1013 vssd1 vssd1 vccd1
+ vccd1 _02290_ sky130_fd_sc_hd__a21o_1
Xhold411 _01220_ vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold422 core.register_file.registers_state\[519\] vssd1 vssd1 vccd1 vccd1 net1741
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10022__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold433 core.register_file.registers_state\[191\] vssd1 vssd1 vccd1 vccd1 net1752
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold444 core.register_file.registers_state\[292\] vssd1 vssd1 vccd1 vccd1 net1763
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 core.register_file.registers_state\[537\] vssd1 vssd1 vccd1 vccd1 net1774
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 core.register_file.registers_state\[854\] vssd1 vssd1 vccd1 vccd1 net1785
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 core.register_file.registers_state\[748\] vssd1 vssd1 vccd1 vccd1 net1796
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_2
X_09944_ net2178 core.CPU_DAT_O\[0\] net800 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XANTENNA__06241__A2 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold488 core.register_file.registers_state\[431\] vssd1 vssd1 vccd1 vccd1 net1807
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 _01449_ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_2
Xhold499 core.register_file.registers_state\[806\] vssd1 vssd1 vccd1 vccd1 net1818
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1113_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout924 net925 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__buf_4
XANTENNA__09715__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout935 net936 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_2
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08140__A _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _04957_ net384 net266 net2138 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__a22o_1
Xfanout957 _01374_ vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10325__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout968 _01372_ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_5_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 core.register_file.registers_state\[351\] vssd1 vssd1 vccd1 vccd1 net2419
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 net981 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_2
Xhold1111 core.register_file.registers_state\[848\] vssd1 vssd1 vccd1 vccd1 net2430
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 core.register_file.registers_state\[168\] vssd1 vssd1 vccd1 vccd1 net2441
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net567 _04711_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__and3_1
Xhold1133 core.register_file.registers_state\[23\] vssd1 vssd1 vccd1 vccd1 net2452
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 core.register_file.registers_state\[667\] vssd1 vssd1 vccd1 vccd1 net2463
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 core.register_file.registers_state\[734\] vssd1 vssd1 vccd1 vccd1 net2474
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 core.register_file.registers_state\[859\] vssd1 vssd1 vccd1 vccd1 net2485
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_120_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ core.IO_mod.input_reg\[19\] net252 net725 vssd1 vssd1 vccd1 vccd1 _04813_
+ sky130_fd_sc_hd__a21o_1
Xhold1177 _01215_ vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
X_05969_ _02067_ _02068_ _02069_ net651 net1004 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a221o_1
Xhold1188 core.register_file.registers_state\[323\] vssd1 vssd1 vccd1 vccd1 net2507
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_A _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 core.register_file.registers_state\[212\] vssd1 vssd1 vccd1 vccd1 net2518
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ _03543_ _03812_ _03480_ _03510_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_105_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ core.IO_mod.data_from_mem\[8\] net249 _04754_ vssd1 vssd1 vccd1 vccd1 _04755_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09494__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ net452 _02931_ net444 net509 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10650_ clknet_leaf_5_clk _00162_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_118_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09246__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09309_ _04931_ net417 net332 net1924 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ clknet_leaf_62_clk _00093_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06480__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08757__A1 core.IO_mod.input_reg\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ clknet_leaf_78_clk _00714_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06217__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11133_ clknet_leaf_19_clk _00645_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[605\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05674__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ clknet_leaf_10_clk _00576_ net1149 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[536\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05991__A1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ net594 _01925_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__nor2_1
XANTENNA__07193__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06091__S1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09485__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917_ clknet_leaf_100_clk _00429_ net1165 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[389\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07496__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07496__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10848_ clknet_leaf_52_clk _00360_ net1304 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[320\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10779_ clknet_leaf_25_clk _00291_ net1186 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08996__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout209 _04334_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_07990_ _03688_ _04084_ _04089_ _04025_ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09056__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ core.register_file.registers_state\[555\] core.register_file.registers_state\[523\]
+ net833 vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05982__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05982__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ _04786_ net286 net282 net2284 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__a22o_1
X_06872_ net1088 _02975_ _02976_ net1067 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ _04004_ _04043_ _04287_ _04298_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nand4_1
XANTENNA__07723__A2 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05823_ net1090 net897 _01867_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a21o_1
XANTENNA__05734__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ _04947_ net395 net299 net1901 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05734__B2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ _01584_ _04612_ _04616_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10857__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05754_ net1032 _01857_ _01858_ _01854_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__o22a_1
XANTENNA__11490__SET_B net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06619__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09476__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ core.pc.current_pc\[22\] _04540_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__and2_1
XANTENNA__09997__Y _05099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05750__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05685_ net949 core.register_file.registers_state\[629\] net763 _01789_ vssd1 vssd1
+ vccd1 vccd1 _01790_ sky130_fd_sc_hd__o31a_1
XFILLER_0_134_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05498__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06695__C1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ net816 _03525_ _03524_ net784 vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09228__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10726__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07239__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07355_ _03453_ _03454_ net1083 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout321_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1063_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05759__A _01862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08987__A1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06306_ net1031 _02408_ _02410_ net1006 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07286_ _03260_ _03263_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06998__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09025_ net745 net464 _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06237_ net633 _02340_ _02341_ net719 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__a211o_1
XANTENNA__06462__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout207_X net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1230_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09936__A0 core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05670__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 net145 vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08422__X _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06168_ net719 _02271_ _02259_ _02251_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a2bb2o_2
Xhold241 net175 vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 net152 vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 _01207_ vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 net190 vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06214__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold285 core.register_file.registers_state\[260\] vssd1 vssd1 vccd1 vccd1 net1604
+ sky130_fd_sc_hd__dlygate4sd3_1
X_06099_ net717 _02182_ _02190_ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__o31a_4
Xhold296 core.register_file.registers_state\[653\] vssd1 vssd1 vccd1 vccd1 net1615
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1116_X net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_33_clk_X clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout721 net722 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_8
XANTENNA__05422__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07962__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 _01419_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
X_09927_ net1082 core.CPU_DAT_O\[16\] net891 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XANTENNA__05973__A1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout743 net745 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_4
XANTENNA_fanout955_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_4
Xfanout776 _01463_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
X_09858_ _04923_ net385 net266 net2032 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__a22o_1
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout798 net801 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06102__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07175__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08809_ net1952 net466 net432 _04857_ vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ _04765_ net385 net273 net2078 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ clknet_leaf_54_clk _01321_ net1299 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09467__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11751_ clknet_leaf_32_clk _01263_ net1206 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
X_10702_ clknet_leaf_89_clk _00214_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[174\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06686__C1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11682_ clknet_leaf_32_clk _01194_ net1205 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06150__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05584__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09219__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10633_ clknet_leaf_38_clk _00145_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07868__B _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_106_clk_X clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07325__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10564_ clknet_leaf_77_clk _00076_ net1261 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10495_ net1413 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09927__A0 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07089__S0 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07402__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ clknet_leaf_105_clk _00628_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[588\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11047_ clknet_leaf_90_clk _00559_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[519\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09604__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05716__A1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06439__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_71_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08130__A2 _03890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05470_ net616 _01573_ _01574_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ net994 core.register_file.registers_state\[452\] net884 core.register_file.registers_state\[484\]
+ net983 vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11505__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09091__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05298__B core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07071_ _03172_ _03174_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10240__A3 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05878__S1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09918__A0 core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__A _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06022_ _02123_ _02124_ _02126_ _02125_ net636 net620 vssd1 vssd1 vccd1 vccd1 _02127_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06902__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08197__A2 _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07973_ _03775_ _03778_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05955__A1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09712_ _05026_ _05062_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__or2_4
X_06924_ core.register_file.registers_state\[43\] net832 vssd1 vssd1 vccd1 vccd1 _03029_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07157__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ net999 _05019_ net461 net393 net1903 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__a32o_1
X_06855_ _02956_ _02957_ _02959_ _02958_ net792 net827 vssd1 vssd1 vccd1 vccd1 _02960_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout271_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A _04898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05806_ net1060 core.register_file.registers_state\[178\] net690 core.register_file.registers_state\[146\]
+ net649 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a221o_1
X_09574_ _04913_ net401 net300 net2239 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06786_ net1097 core.register_file.registers_state\[976\] core.register_file.registers_state\[1008\]
+ net839 net1073 vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__o221a_1
XANTENNA__09449__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06380__B2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08525_ _04588_ _04597_ _04599_ _04596_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a31o_1
XANTENNA__11035__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05737_ net662 _01840_ _01841_ net965 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06668__C1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1278_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08456_ _04540_ _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__nor2_1
X_05668_ net1057 core.register_file.registers_state\[470\] vssd1 vssd1 vccd1 vccd1
+ _01773_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06132__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06132__B2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07407_ _03509_ _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__nand2_1
XANTENNA__08409__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ core.pc.current_pc\[14\] _04479_ net599 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__mux2_1
XANTENNA__07880__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05599_ net638 _01700_ _01701_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout703_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_X net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07338_ net1095 core.register_file.registers_state\[859\] core.register_file.registers_state\[891\]
+ net836 net979 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__o221a_1
XANTENNA__09082__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09621__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07093__C1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07269_ net778 _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09909__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ net2517 net428 _04978_ net434 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__a22o_1
XANTENNA__06840__C1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ net33 net903 net795 net2068 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10334__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__B _04401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07991__X _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05655__C net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_2
Xfanout562 _04712_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
Xfanout573 _04668_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_4
Xfanout584 _01505_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_13_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_2
XFILLER_0_9_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09143__B net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10648__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11803_ clknet_leaf_70_clk _01304_ net1275 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_53_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08982__B _04662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ clknet_leaf_46_clk _01246_ net1289 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11528__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09860__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ clknet_leaf_45_clk _01177_ net1289 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07598__B _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10616_ clknet_leaf_5_clk _00128_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ clknet_leaf_27_clk _01108_ net1203 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09612__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10552__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10547_ clknet_leaf_97_clk _00059_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10222__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10478_ net1400 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08179__A2 _03959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07387__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A2 _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05937__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09037__C _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07139__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11058__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09053__B _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ net778 _02738_ _02739_ net773 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a31o_1
XANTENNA__06362__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10199__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06396__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06571_ net1095 core.register_file.registers_state\[87\] core.register_file.registers_state\[119\]
+ net836 net803 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__o221a_1
XANTENNA__05570__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08310_ _02207_ _04407_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05522_ _01399_ _01500_ _01614_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__or3_1
X_09290_ net2514 net243 net336 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06114__A1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09851__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05801__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08241_ core.pc.current_pc\[0\] net575 vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__nor2_1
X_05453_ net1043 core.register_file.registers_state\[733\] core.register_file.registers_state\[765\]
+ net672 net653 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08172_ _03774_ _03889_ _03909_ _03798_ _04276_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__o221a_1
X_05384_ net1003 net896 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__nor2_4
XFILLER_0_16_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09603__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07123_ _03226_ _03227_ net974 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07728__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06822__C1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ net974 _03155_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__a21o_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_11_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06005_ net1013 _02107_ _02108_ net963 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09367__B2 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_112_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1026_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_11_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__07029__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput198 net198 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__05928__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout486_A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _03826_ _04018_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07316__X _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06907_ core.register_file.registers_state\[12\] core.register_file.registers_state\[44\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07887_ _03821_ _03925_ _03969_ _03991_ net479 net495 vssd1 vssd1 vccd1 vccd1 _03992_
+ sky130_fd_sc_hd__mux4_2
XANTENNA_fanout653_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06838_ core.register_file.registers_state\[47\] core.register_file.registers_state\[15\]
+ net848 vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
X_09626_ net744 _04997_ net460 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09557_ net205 net2477 net303 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06769_ _01987_ _02842_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout820_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08508_ _04585_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06807__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06105__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09488_ net603 _04892_ net316 net261 net1908 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_82_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08439_ _01896_ _04511_ _04515_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10329__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07853__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05864__B1 core.register_file.registers_state\[369\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ clknet_leaf_7_clk _00962_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_134_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ net1419 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_134_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10204__A3 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08802__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ clknet_leaf_63_clk _00893_ net1249 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10332_ _05117_ net1593 net240 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08323__A core.decoder.inst\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10263_ net2252 _05239_ _04360_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07369__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1302 net1305 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__clkbuf_4
X_10194_ net122 net918 net909 net1595 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__a22o_1
XANTENNA__08030__B2 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A gpio_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05919__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06041__A0 _02117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1313 net1314 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__buf_4
XFILLER_0_100_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08977__B net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 _04898_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_2
XANTENNA__06592__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout381 net382 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_6
XANTENNA__05682__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout392 _05066_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08604__D_N _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10918__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09294__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ clknet_leaf_50_clk net1500 net1308 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07844__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11648_ clknet_leaf_50_clk _01160_ net1307 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_2
XFILLER_0_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07057__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput45 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11579_ clknet_leaf_29_clk _01091_ net1200 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[27\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput56 gpio_in[29] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput67 nrst vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_1
Xhold807 core.register_file.registers_state\[109\] vssd1 vssd1 vccd1 vccd1 net2126
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold818 core.register_file.registers_state\[480\] vssd1 vssd1 vccd1 vccd1 net2137
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11270__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold829 core.register_file.registers_state\[122\] vssd1 vssd1 vccd1 vccd1 net2148
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09349__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09048__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08557__C1 _01508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06258__S1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ _03697_ _03891_ _03905_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__o211a_2
X_08790_ net727 _03916_ net525 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__a21o_1
XANTENNA__06583__A1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06688__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__C_N _04317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _02519_ _03662_ _03663_ _03797_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09064__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06040__X _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A1 _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ net452 _02962_ net444 net506 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09999__A _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__X _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ net2220 net206 net406 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
XANTENNA__10598__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06623_ core.register_file.registers_state\[917\] core.register_file.registers_state\[949\]
+ net879 vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11843__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ _04982_ net416 net412 net1624 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a22o_1
XANTENNA__08088__A1 _03622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06554_ net769 _02658_ _02646_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05505_ net934 _01606_ _01609_ net719 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a31o_1
XANTENNA__07835__A1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ net2500 _04890_ net335 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__mux2_1
X_06485_ _02586_ _02589_ net631 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout234_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09938__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08224_ _01628_ _03742_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05436_ net617 _01539_ _01540_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__or3_1
XANTENNA__08842__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07048__C1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08155_ _02935_ _04005_ _02998_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o21ai_1
X_05367_ net1099 core.register_file.registers_state\[478\] core.register_file.registers_state\[510\]
+ net841 net1073 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout401_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1143_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07106_ net1098 core.register_file.registers_state\[677\] core.register_file.registers_state\[645\]
+ net842 net805 vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08260__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ net1113 _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nor2_1
X_05298_ core.decoder.inst\[25\] core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1 _01413_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_101_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11223__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07037_ _03139_ _03141_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1029_X net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06598__A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net614 net225 vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__and2_1
XANTENNA__06574__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07939_ _03397_ _03399_ _03144_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05933__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05782__C1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09512__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ clknet_leaf_99_clk _00462_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[422\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ _04974_ net397 net392 net1936 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ clknet_leaf_86_clk _00393_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[353\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07826__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11502_ clknet_leaf_66_clk _01014_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[974\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11433_ clknet_leaf_17_clk _00945_ net1211 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[905\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10189__A2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11467__SET_B net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11364_ clknet_leaf_81_clk _00876_ net1255 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[836\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08053__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06262__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10315_ _05100_ net1529 net237 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11295_ clknet_leaf_16_clk _00807_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[767\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08988__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10246_ net1126 net1437 net911 _05231_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__a31o_1
XANTENNA__08003__A1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1110 core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_4
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_2
Xfanout1132 net1134 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_4
X_10177_ net104 net916 net906 net1465 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a22o_1
Xfanout1143 net1145 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__clkbuf_4
Xfanout1154 net1157 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06565__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_2
Xfanout1176 net1177 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
Xfanout1187 net1209 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05773__C1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1198 net1202 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09503__A1 _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06317__A1 _01506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__X _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06270_ net1059 core.register_file.registers_state\[484\] net754 _02374_ vssd1 vssd1
+ vccd1 vccd1 _02375_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07045__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold604 core.register_file.registers_state\[520\] vssd1 vssd1 vccd1 vccd1 net1923
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09059__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold615 core.register_file.registers_state\[698\] vssd1 vssd1 vccd1 vccd1 net1934
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 core.register_file.registers_state\[634\] vssd1 vssd1 vccd1 vccd1 net1945
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold637 core.register_file.registers_state\[556\] vssd1 vssd1 vccd1 vccd1 net1956
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 core.register_file.registers_state\[692\] vssd1 vssd1 vccd1 vccd1 net1967
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ core.IO_mod.data_from_mem\[16\] core.CPU_DAT_O\[16\] net799 vssd1 vssd1 vccd1
+ vccd1 _01112_ sky130_fd_sc_hd__mux2_1
Xhold659 net173 vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09990__B2 _02421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ _04758_ net602 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__nor2_1
X_09891_ net1115 _04986_ net457 net375 net1683 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload19_A clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06005__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ net226 net2354 net373 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08773_ _04670_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__nor2_1
X_05985_ core.register_file.registers_state\[524\] core.register_file.registers_state\[556\]
+ net698 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
XANTENNA__05764__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ net1003 _01708_ _03446_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10104__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ net506 net449 _03351_ net441 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__or4_1
XANTENNA__06403__S1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1093_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06606_ net783 _02709_ _02710_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__or3_1
X_07586_ _01501_ _01626_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__or2_1
XANTENNA__09258__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__A _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ _04955_ net420 net333 net2088 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06537_ net1104 core.register_file.registers_state\[348\] core.register_file.registers_state\[380\]
+ net850 net982 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__o221a_1
XFILLER_0_36_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11560__Q core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout616_A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05819__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ net560 _04877_ _05044_ net341 net2087 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06468_ _02565_ _02571_ _02572_ _02564_ net932 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08207_ _01393_ _01395_ _01868_ net546 _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05419_ net1029 net753 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__nand2_4
XFILLER_0_90_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09187_ _04979_ net355 net424 net2480 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06399_ net946 core.register_file.registers_state\[65\] net702 core.register_file.registers_state\[97\]
+ net657 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08138_ _04229_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout985_A _01370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10040__B2 _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08069_ _03392_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1313_X net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10100_ net1452 net516 _05159_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11080_ clknet_leaf_12_clk _00592_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[552\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_129_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08601__A _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net724 _01646_ _01663_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__and3_4
XANTENNA__10342__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11119__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ clknet_leaf_62_clk _00445_ net1242 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[405\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10864_ clknet_leaf_107_clk _00376_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[336\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09249__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10795_ clknet_leaf_108_clk _00307_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08054__Y _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11416_ clknet_leaf_4_clk _00928_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[888\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11347_ clknet_leaf_11_clk _00859_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08775__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07983__A0 _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11278_ clknet_leaf_89_clk _00790_ net1235 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[750\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08527__A2 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10229_ net75 net920 vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__and2_1
XANTENNA__06538__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B1 _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06538__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07127__A _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1 core.register_file.registers_state\[938\] vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05746__C1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05770_ net622 _01871_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09488__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07499__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08229__Y _04334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ _03450_ _03478_ _03481_ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_18_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07371_ _03475_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ _04654_ net604 _04714_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__or3_4
X_06322_ net662 _02425_ _02426_ net965 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__o211a_1
XANTENNA__10636__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__X _04350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06905__S net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09660__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09041_ net998 net462 _05000_ net427 net1968 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__a32o_1
X_06253_ net964 _02353_ _02355_ _02357_ net934 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06184_ core.register_file.registers_state\[294\] core.register_file.registers_state\[262\]
+ core.register_file.registers_state\[422\] core.register_file.registers_state\[390\]
+ net674 net1014 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux4_1
Xhold401 core.register_file.registers_state\[542\] vssd1 vssd1 vccd1 vccd1 net1720
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold412 core.register_file.registers_state\[413\] vssd1 vssd1 vccd1 vccd1 net1731
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10786__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06226__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold423 core.register_file.registers_state\[405\] vssd1 vssd1 vccd1 vccd1 net1742
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 net191 vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10022__B2 _05111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold445 core.register_file.registers_state\[404\] vssd1 vssd1 vccd1 vccd1 net1764
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold456 core.register_file.registers_state\[784\] vssd1 vssd1 vccd1 vccd1 net1775
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold467 core.register_file.registers_state\[258\] vssd1 vssd1 vccd1 vccd1 net1786
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold478 core.register_file.registers_state\[774\] vssd1 vssd1 vccd1 vccd1 net1797
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ core.ru.state\[4\] _01441_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__and2_1
Xhold489 core.register_file.registers_state\[816\] vssd1 vssd1 vccd1 vccd1 net1808
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout903 _05243_ vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout936 net943 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout399_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09874_ _04955_ net390 net268 net2106 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__a22o_1
Xfanout947 net957 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 net961 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
XANTENNA__09951__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1106_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 core.register_file.registers_state\[132\] vssd1 vssd1 vccd1 vccd1 net2420
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_4
XANTENNA__07037__A _03139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 core.register_file.registers_state\[605\] vssd1 vssd1 vccd1 vccd1 net2431
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1123 core.register_file.registers_state\[307\] vssd1 vssd1 vccd1 vccd1 net2442
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ net605 _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_2
Xhold1134 core.register_file.registers_state\[316\] vssd1 vssd1 vccd1 vccd1 net2453
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1145 core.register_file.registers_state\[595\] vssd1 vssd1 vccd1 vccd1 net2464
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 core.register_file.registers_state\[660\] vssd1 vssd1 vccd1 vccd1 net2475
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 core.register_file.registers_state\[604\] vssd1 vssd1 vccd1 vccd1 net2486
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05968_ net923 _02070_ _02072_ net932 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a211o_1
Xhold1178 core.register_file.registers_state\[658\] vssd1 vssd1 vccd1 vccd1 net2497
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ net2152 net469 net439 _04812_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_120_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 core.register_file.registers_state\[592\] vssd1 vssd1 vccd1 vccd1 net2508
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09252__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07707_ _03421_ _03422_ _03540_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08687_ core.IO_mod.input_reg\[8\] net253 net730 vssd1 vssd1 vccd1 vccd1 _04754_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_105_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05899_ net951 core.register_file.registers_state\[847\] net709 core.register_file.registers_state\[879\]
+ net1020 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09494__A3 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07638_ _02606_ _03549_ net527 vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06087__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06162__C1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06701__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06701__B2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ net455 _03506_ net447 vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09308_ _04929_ net419 net333 net1997 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10580_ clknet_leaf_55_clk _00092_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09651__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ net560 _04834_ _05035_ net341 net2396 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08315__B _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06560__S0 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ clknet_leaf_85_clk _00713_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[673\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06217__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__A1 _01978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06768__A1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ clknet_leaf_42_clk _00644_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[604\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold990 core.register_file.registers_state\[141\] vssd1 vssd1 vccd1 vccd1 net2309
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05440__B2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ clknet_leaf_21_clk _00575_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[535\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10014_ net1533 net542 net521 _05107_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09182__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07193__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__B net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07732__A3 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06940__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05743__A2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10659__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__A_N _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10916_ clknet_leaf_80_clk _00428_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[388\]
+ sky130_fd_sc_hd__dfrtp_1
X_11896_ net136 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09890__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05900__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10847_ clknet_leaf_14_clk _00359_ net1175 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[319\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10778_ clknet_leaf_7_clk _00290_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[250\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09642__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10252__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08996__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10004__B2 _05102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06940_ net970 _03041_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__a21o_1
XANTENNA__09056__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09173__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06871_ net991 core.register_file.registers_state\[718\] net878 core.register_file.registers_state\[750\]
+ net808 vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11884__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11434__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__B2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _03884_ _04684_ _03985_ _03862_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__or4bb_1
X_05822_ net1087 net897 _01867_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a21oi_2
X_09590_ _04945_ net396 net299 net2242 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__a22o_1
XANTENNA__08387__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09072__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ core.pc.current_pc\[28\] net595 _04617_ _04619_ vssd1 vssd1 vccd1 vccd1 _00036_
+ sky130_fd_sc_hd__o22a_1
X_05753_ net1023 _01855_ _01856_ net965 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08472_ _04553_ _04555_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11584__CLK clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06144__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__A _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05684_ net1054 core.register_file.registers_state\[597\] vssd1 vssd1 vccd1 vccd1
+ _01789_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09881__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05498__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload86_A clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07423_ _03526_ _03527_ net791 vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07354_ _03455_ _03456_ _03457_ _03458_ net784 net803 vssd1 vssd1 vccd1 vccd1 _03459_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08416__A _01958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06305_ net1062 core.register_file.registers_state\[739\] net755 _02409_ net929 vssd1
+ vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a311o_1
XANTENNA__06447__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08987__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ _03387_ _03388_ _03293_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout314_A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06998__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06542__S0 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1056_A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ net613 net220 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__and2_1
XANTENNA__09946__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06236_ net622 _02333_ _02334_ _02331_ net627 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__o311a_1
XFILLER_0_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08168__A1_N net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold220 core.register_file.registers_state\[0\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06167_ _02251_ _02259_ _02271_ net719 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__o2bb2a_2
Xhold231 core.ADR_I\[4\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 core.register_file.registers_state\[926\] vssd1 vssd1 vccd1 vccd1 net1561
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 core.CPU_DAT_I\[20\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 core.IO_mod.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08151__A _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 core.IO_mod.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
X_06098_ net632 _02195_ _02202_ net717 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__o211ai_1
XANTENNA__05958__C1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold286 core.register_file.registers_state\[551\] vssd1 vssd1 vccd1 vccd1 net1605
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_4
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05422__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 core.register_file.registers_state\[406\] vssd1 vssd1 vccd1 vccd1 net1616
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 net715 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07962__A3 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09926_ net1095 net2555 net891 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
Xfanout722 _01511_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_6
Xfanout733 _01419_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1109_X net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout755 net756 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_4
XANTENNA__09164__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 _01509_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_4
XANTENNA_fanout850_A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _04921_ net383 net266 net1658 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__a22o_1
Xfanout777 net778 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout788 _01456_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
XANTENNA__07175__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout799 net801 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08808_ net565 _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _04760_ net385 net270 net1823 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ core.IO_mod.input_reg\[16\] net250 net725 vssd1 vssd1 vccd1 vccd1 _04798_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ clknet_leaf_32_clk _01262_ net1206 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09872__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ clknet_leaf_2_clk _00213_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[173\]
+ sky130_fd_sc_hd__dfrtp_1
X_11681_ clknet_leaf_32_clk _01193_ net1207 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05584__S1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10632_ clknet_leaf_14_clk _00144_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10234__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10563_ clknet_leaf_73_clk _00075_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08045__B _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05388__C core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10494_ net1376 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07089__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07938__B1 _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07402__A2 _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06205__A3 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__B_N _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05949__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05413__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ clknet_leaf_107_clk _00627_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[587\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06610__B1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05413__B2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09155__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11046_ clknet_leaf_99_clk _00558_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[518\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10170__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06913__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06913__B2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11224__RESET_B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07899__X _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09863__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11879_ clknet_leaf_71_clk _01348_ net1276 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06772__S0 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06429__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07070_ _03172_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06021_ core.register_file.registers_state\[1003\] core.register_file.registers_state\[971\]
+ net667 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__B _03536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09067__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05404__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07972_ _03657_ _03951_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05882__X _01987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ net241 net2172 net281 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
X_06923_ net1092 core.register_file.registers_state\[139\] net832 core.register_file.registers_state\[171\]
+ net816 vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__o221a_1
XANTENNA__07157__A1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09642_ _05017_ net396 net391 net2335 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__a22o_1
X_06854_ core.register_file.registers_state\[943\] core.register_file.registers_state\[911\]
+ net853 vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__mux2_1
X_05805_ net1007 _01900_ _01904_ _01909_ net630 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_102_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06785_ net1097 core.register_file.registers_state\[848\] core.register_file.registers_state\[880\]
+ net839 net980 vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__o221a_1
X_09573_ _04911_ net397 net302 net1941 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout264_A _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08524_ core.pc.current_pc\[27\] _04592_ net228 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__o21ai_1
X_05736_ net1063 core.register_file.registers_state\[724\] vssd1 vssd1 vccd1 vccd1
+ _01841_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08845__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09854__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08455_ core.pc.current_pc\[20\] _04520_ core.pc.current_pc\[21\] vssd1 vssd1 vccd1
+ vccd1 _04541_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05667_ net949 core.register_file.registers_state\[374\] net764 _01771_ net928 vssd1
+ vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout431_A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1173_A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07406_ _03506_ _03508_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__nand2_1
X_08386_ _04478_ _04477_ _04476_ net209 vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_107_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05598_ net937 core.register_file.registers_state\[251\] net748 _01702_ net1010 vssd1
+ vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10216__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07337_ net1095 core.register_file.registers_state\[987\] core.register_file.registers_state\[1019\]
+ net837 net1071 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ net977 _03369_ _03372_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06219_ core.register_file.registers_state\[293\] core.register_file.registers_state\[261\]
+ core.register_file.registers_state\[421\] core.register_file.registers_state\[389\]
+ net682 net1017 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux4_1
XANTENNA__09909__A1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ net565 _04977_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07199_ net976 _03294_ _03303_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1226_X net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09385__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout530 _03624_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_4
Xfanout541 net543 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_2
X_09909_ net1117 _05019_ net461 net377 net1561 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__a32o_1
Xfanout563 net566 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_4
Xfanout574 _04336_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08345__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 net587 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
Xfanout596 net600 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10350__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__B1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06356__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11802_ clknet_leaf_71_clk _01303_ net1271 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ clknet_leaf_45_clk _01245_ net1289 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07320__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07320__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11664_ clknet_leaf_45_clk _01176_ net1289 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05882__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ clknet_leaf_22_clk _00127_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11595_ clknet_leaf_27_clk _01107_ net1204 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10546_ clknet_leaf_71_clk _00058_ net1274 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output183_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10477_ net1371 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10847__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09376__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06304__A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07926__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07139__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10997__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ clknet_leaf_62_clk _00541_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[501\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10143__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06570_ core.register_file.registers_state\[23\] core.register_file.registers_state\[55\]
+ core.register_file.registers_state\[151\] core.register_file.registers_state\[183\]
+ net866 net818 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09836__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05521_ net1114 _01499_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09300__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08240_ _03351_ _04335_ _04342_ _02488_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05452_ net1043 core.register_file.registers_state\[605\] core.register_file.registers_state\[637\]
+ net672 net638 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05873__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _03890_ _03981_ _04273_ _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11622__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05383_ _01475_ _01487_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__nand2_8
XFILLER_0_16_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07122_ net990 core.register_file.registers_state\[453\] net876 core.register_file.registers_state\[485\]
+ net982 vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload49_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07053_ net1086 _03156_ _03157_ net777 vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_101_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06004_ core.register_file.registers_state\[268\] core.register_file.registers_state\[300\]
+ core.register_file.registers_state\[396\] core.register_file.registers_state\[428\]
+ net698 net1013 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__09367__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_11_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XANTENNA__10007__Y _05104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07378__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XANTENNA__07378__B2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_11_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput199 net199 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1019_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ net490 _04059_ _04054_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout381_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_X clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06906_ net1098 core.register_file.registers_state\[172\] net841 core.register_file.registers_state\[140\]
+ net806 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__a221o_1
XANTENNA__10023__X _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ net502 _03640_ _03647_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09625_ net2505 net394 _05074_ net1000 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11563__Q core.decoder.inst\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ net975 _02938_ _02941_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _04832_ net2386 net304 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__mux2_1
XANTENNA__11152__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09827__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06768_ net774 _02872_ _02861_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a21o_4
XFILLER_0_78_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08507_ _04587_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__nand2b_1
X_05719_ _01811_ _01823_ _01805_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout813_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ core.register_file.registers_state\[275\] core.register_file.registers_state\[307\]
+ core.register_file.registers_state\[403\] core.register_file.registers_state\[435\]
+ net871 net1074 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux4_1
XANTENNA__06105__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _05005_ net322 net264 net1828 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08438_ _04524_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__nand2_1
XANTENNA__07853__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06510__C1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05864__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05864__B2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ core.pc.current_pc\[13\] _02931_ net576 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire227 _04719_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09055__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10400_ net1397 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07066__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11380_ clknet_leaf_57_clk _00892_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[852\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07605__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08604__A _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08802__B2 _04851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10331_ _05116_ net1700 net237 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10345__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08323__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10262_ _04346_ _04347_ _02424_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09358__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07369__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10193_ net121 net919 net909 net1499 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1303 net1304 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06577__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1314 net67 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__buf_6
XANTENNA__05919__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06041__A1 _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06411__X _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout371 _04883_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_89_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout382 _05087_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout393 _05066_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_31_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09530__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ clknet_leaf_46_clk net1546 net1290 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11647_ clknet_leaf_46_clk _01159_ net1290 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07829__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09597__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07057__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11795__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput35 gpio_in[0] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11578_ clknet_leaf_33_clk _01090_ net1203 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[26\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput46 gpio_in[1] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
Xinput57 gpio_in[2] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xhold808 core.register_file.registers_state\[896\] vssd1 vssd1 vccd1 vccd1 net2127
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold819 core.register_file.registers_state\[893\] vssd1 vssd1 vccd1 vccd1 net2138
+ sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ clknet_leaf_84_clk _00041_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08233__B _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06280__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11025__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08801__X _04851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10364__A0 _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08887__C net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06583__A2 _01781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07740_ _03645_ _03646_ _03674_ _03675_ net499 net476 vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09064__B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10116__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05791__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_74_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ net506 _03632_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a21boi_1
XANTENNA__09999__B _02174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__B _02113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ net2304 net222 net405 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
X_06622_ core.register_file.registers_state\[981\] core.register_file.registers_state\[1013\]
+ net879 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XANTENNA__05543__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09809__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__RESET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06553_ net967 _02654_ _02657_ _02651_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a31o_1
X_09341_ _04980_ net418 net413 net1844 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09285__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06099__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_89_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05504_ net645 _01607_ _01608_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ net2257 net206 net336 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__mux2_1
X_06484_ net616 _02587_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__or3_1
XANTENNA__07835__A2 _03939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06209__A _02296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08223_ _04325_ _04326_ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__nor3_1
X_05435_ net1048 core.register_file.registers_state\[222\] core.register_file.registers_state\[254\]
+ net676 net655 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07048__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _04075_ _04109_ _04123_ _04258_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_16_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05366_ net1098 core.register_file.registers_state\[350\] core.register_file.registers_state\[382\]
+ net842 net980 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10198__A3 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07105_ core.register_file.registers_state\[549\] core.register_file.registers_state\[517\]
+ net841 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__mux2_1
XANTENNA__08796__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ net533 _03290_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__or2_1
X_05297_ _01409_ _01411_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__or2_4
XANTENNA__09954__S net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07036_ _02241_ _03112_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11558__Q core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10355__A0 _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1303_A net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06559__C1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09760__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ net1002 net464 _04964_ net429 net2122 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A1 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10107__B1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07938_ _04029_ _04030_ _04039_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_127_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10542__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11668__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07869_ net532 _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a21boi_1
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08720__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ _04972_ net399 net392 net2067 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10880_ clknet_leaf_51_clk _00392_ net1304 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[352\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06818__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05534__B1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07503__A _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09539_ _04884_ net2281 net305 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09276__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11501_ clknet_leaf_0_clk _01013_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[973\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_109_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09579__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ clknet_leaf_9_clk _00944_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11363_ clknet_leaf_65_clk _00875_ net1245 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[835\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ _05099_ net1642 net238 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11294_ clknet_leaf_95_clk _00806_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08988__B net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ net84 net914 vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10346__A0 _05098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1102 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05693__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07211__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1111 core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_4
Xfanout1122 core.decoder.inst\[9\] vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09751__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ net103 net916 net906 net1667 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__a22o_1
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_4
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07762__A1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1155 net1157 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
Xfanout1166 net1167 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_2
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_2
Xfanout1188 net1190 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__clkbuf_4
Xfanout1199 net1202 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05980__X _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06970__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09503__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06317__A2 _02421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload5_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09267__A1 _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09806__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09059__B _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold605 core.register_file.registers_state\[368\] vssd1 vssd1 vccd1 vccd1 net1924
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06789__C1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold616 core.register_file.registers_state\[649\] vssd1 vssd1 vccd1 vccd1 net1935
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold627 core.register_file.registers_state\[153\] vssd1 vssd1 vccd1 vccd1 net1946
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 core.register_file.registers_state\[60\] vssd1 vssd1 vccd1 vccd1 net1957
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06253__A1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold649 core.register_file.registers_state\[147\] vssd1 vssd1 vccd1 vccd1 net1968
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11420__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09990__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ net2313 net369 _04913_ net437 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__a22o_1
X_09890_ net1115 _05070_ net375 net2415 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__a22o_1
XANTENNA__06005__A1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09075__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ net207 net2367 net374 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__mux2_1
XANTENNA__09742__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07753__B2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ _04823_ _04824_ _04825_ _04757_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__a211o_2
X_05984_ core.register_file.registers_state\[780\] core.register_file.registers_state\[812\]
+ core.register_file.registers_state\[908\] core.register_file.registers_state\[940\]
+ net697 net1014 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux4_1
XANTENNA__05764__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ _01708_ _03446_ net580 vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07654_ net494 _03757_ _03751_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06713__C1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06605_ net825 _02706_ _02705_ net786 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11473__SET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09258__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ net265 _03689_ _03682_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout344_A _05027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__B _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1086_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09949__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _04953_ net418 net331 net2347 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06536_ core.register_file.registers_state\[284\] core.register_file.registers_state\[316\]
+ core.register_file.registers_state\[412\] core.register_file.registers_state\[444\]
+ net881 net1077 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux4_1
XANTENNA__08853__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ core.register_file.registers_state\[318\] net475 net545 vssd1 vssd1 vccd1
+ vccd1 _05044_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout511_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06467_ net936 core.register_file.registers_state\[824\] net760 net923 vssd1 vssd1
+ vccd1 vccd1 _02572_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout1253_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout609_A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _01895_ net550 vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05418_ net960 net761 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__nor2_1
X_06398_ _02500_ _02502_ net618 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09186_ _04977_ net355 net424 net1963 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05349_ core.i_hit _01437_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_116_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08137_ _04022_ _04241_ _04240_ _04235_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__o211a_4
XFILLER_0_47_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09430__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11340__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_X net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10040__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08068_ _03234_ _03235_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout880_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05452__C1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__A0 _05113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07019_ net972 _03122_ _03123_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_129_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10030_ net1779 net543 net522 _05115_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__a22o_1
XANTENNA__09194__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09733__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05755__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05507__A0 _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ clknet_leaf_55_clk _00444_ net1295 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[404\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06704__C1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11751__Q net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ clknet_leaf_84_clk _00375_ net1232 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[335\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09249__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08616__X _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10794_ clknet_leaf_106_clk _00306_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08209__C1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06483__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06483__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ clknet_leaf_22_clk _00927_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[887\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09421__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08214__D _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ clknet_leaf_67_clk _00858_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[818\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11833__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__A0 _05104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11277_ clknet_leaf_3_clk _00789_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09185__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10228_ net1127 net1424 net912 _05222_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__a31o_1
XANTENNA__09724__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__C1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10884__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07127__B _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10159_ _01450_ _01453_ _05204_ core.BUSY_O vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__o22a_1
Xhold2 core.register_file.registers_state\[954\] vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10813__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06943__C1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09488__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08160__A1 _03791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11546__SET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07370_ _03467_ _03474_ net767 _03462_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_128_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06321_ net1065 core.register_file.registers_state\[672\] core.register_file.registers_state\[640\]
+ net692 net648 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06252_ net660 _02348_ _02356_ net1031 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__a31o_1
X_09040_ net746 net612 net215 vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__and3_1
XANTENNA__11363__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06183_ _02287_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10009__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold402 core.register_file.registers_state\[288\] vssd1 vssd1 vccd1 vccd1 net1721
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 core.register_file.registers_state\[306\] vssd1 vssd1 vccd1 vccd1 net1732
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10022__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold424 net119 vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold435 core.register_file.registers_state\[298\] vssd1 vssd1 vccd1 vccd1 net1754
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold446 core.register_file.registers_state\[271\] vssd1 vssd1 vccd1 vccd1 net1765
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold457 core.register_file.registers_state\[563\] vssd1 vssd1 vccd1 vccd1 net1776
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05434__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold468 core.register_file.registers_state\[297\] vssd1 vssd1 vccd1 vccd1 net1787
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ core.decoder.inst\[31\] core.CPU_DAT_O\[31\] net893 vssd1 vssd1 vccd1 vccd1
+ _01095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold479 core.register_file.registers_state\[696\] vssd1 vssd1 vccd1 vccd1 net1798
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 _05242_ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_2
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout915 net921 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09176__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout926 net931 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09873_ _04953_ net384 net266 net1951 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__a22o_1
Xfanout937 net938 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout948 net949 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07726__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07726__B2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net961 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
X_08824_ net526 _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_5_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 core.register_file.registers_state\[145\] vssd1 vssd1 vccd1 vccd1 net2421
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 core.register_file.registers_state\[640\] vssd1 vssd1 vccd1 vccd1 net2432
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05737__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 core.register_file.registers_state\[68\] vssd1 vssd1 vccd1 vccd1 net2443
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1135 core.register_file.registers_state\[192\] vssd1 vssd1 vccd1 vccd1 net2454
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07752__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1146 core.register_file.registers_state\[680\] vssd1 vssd1 vccd1 vccd1 net2465
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1157 core.register_file.registers_state\[451\] vssd1 vssd1 vccd1 vccd1 net2476
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net571 net609 net216 vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__and3_2
X_05967_ core.register_file.registers_state\[909\] net694 _02071_ vssd1 vssd1 vccd1
+ vccd1 _02072_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout461_A _05060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 core.register_file.registers_state\[499\] vssd1 vssd1 vccd1 vccd1 net2487
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_120_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1179 core.register_file.registers_state\[84\] vssd1 vssd1 vccd1 vccd1 net2498
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _03550_ _03743_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_135_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10031__X _05116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09252__B net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ net1810 net468 net436 _04753_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05898_ net633 _01999_ _02002_ net718 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__o31a_1
X_07637_ _01616_ _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__and2b_1
XANTENNA__11571__Q core.decoder.inst\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout726_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08065__A_N _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_X net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07568_ net498 _03670_ _03672_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06892__A _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09100__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09307_ _04927_ net419 net333 net2057 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06519_ net987 core.register_file.registers_state\[701\] net868 core.register_file.registers_state\[669\]
+ net823 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_118_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07499_ net972 _03600_ _03603_ net776 vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06465__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09238_ core.register_file.registers_state\[310\] _04666_ net545 vssd1 vssd1 vccd1
+ vccd1 _05035_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11342__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05301__A core.decoder.inst\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06560__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09403__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ _04946_ net352 net343 net2033 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06217__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ clknet_leaf_56_clk _00712_ net1286 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[672\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10013__A2 _01985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08612__A _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__A1 _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05425__C1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11131_ clknet_leaf_23_clk _00643_ net1184 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[603\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10353__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 core.register_file.registers_state\[199\] vssd1 vssd1 vccd1 vccd1 net2299
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09167__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold991 core.register_file.registers_state\[718\] vssd1 vssd1 vccd1 vccd1 net2310
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ clknet_leaf_60_clk _00574_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[534\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10013_ _01978_ _01985_ net724 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__o21a_2
XFILLER_0_21_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10915_ clknet_leaf_74_clk _00427_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[387\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11895_ net136 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09890__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10846_ clknet_leaf_92_clk _00358_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[318\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05900__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07102__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10777_ clknet_leaf_54_clk _00289_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[249\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06456__A1 _02560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08081__X _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09618__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10263__S _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ clknet_leaf_85_clk _00841_ net1236 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06042__A core.decoder.inst\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06870_ net992 core.register_file.registers_state\[590\] net878 core.register_file.registers_state\[622\]
+ net824 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__a221o_1
XANTENNA__06977__A _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05881__A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05821_ _01897_ _01925_ net585 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XANTENNA__05814__S0 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08540_ net208 _04618_ net595 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09072__B net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05752_ core.register_file.registers_state\[276\] core.register_file.registers_state\[308\]
+ core.register_file.registers_state\[404\] core.register_file.registers_state\[436\]
+ net714 net1022 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08133__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08471_ _04535_ _04554_ _04553_ _04545_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06144__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05683_ net948 core.register_file.registers_state\[757\] net753 _01787_ net1022 vssd1
+ vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09881__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__B _01956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06695__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07422_ net1091 core.register_file.registers_state\[216\] core.register_file.registers_state\[248\]
+ net835 net816 vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07892__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06695__B2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08256__X _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10753__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07353_ core.register_file.registers_state\[26\] core.register_file.registers_state\[58\]
+ net866 vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11879__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09633__B2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06304_ net955 core.register_file.registers_state\[707\] vssd1 vssd1 vccd1 vccd1
+ _02409_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07284_ _03293_ _03388_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09023_ net2309 net427 _04988_ net431 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__a22o_1
XANTENNA__06542__S1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06235_ _02336_ _02337_ _02338_ _02339_ net625 net643 vssd1 vssd1 vccd1 vccd1 _02340_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1049_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 net172 vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06166_ net934 _02264_ _02267_ _02270_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__o22a_1
Xhold221 core.CPU_DAT_I\[2\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06651__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 net194 vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07947__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold243 net154 vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _01221_ vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 net198 vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
X_06097_ net961 _02196_ _02201_ net628 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a211o_1
Xhold276 core.CPU_DAT_I\[29\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08151__B _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 net195 vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09962__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 net716 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09149__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09925_ core.decoder.inst\[14\] core.CPU_DAT_O\[14\] net892 vssd1 vssd1 vccd1 vccd1
+ _01078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout712 net713 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_4
Xhold298 core.register_file.registers_state\[409\] vssd1 vssd1 vccd1 vccd1 net1617
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout723 _01511_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_6
XANTENNA__11566__Q core.decoder.inst\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11259__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout734 _01412_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout676_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 net746 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_4
Xfanout756 _01510_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_4
Xfanout767 net770 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_6
X_09856_ _04919_ net383 net266 net1757 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 _01463_ vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout789 net791 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07482__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ net605 _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09787_ _04753_ net387 net271 net1736 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout843_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ core.register_file.registers_state\[521\] core.register_file.registers_state\[553\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
X_08738_ net1827 net468 net436 _04797_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09321__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ core.IO_mod.input_reg\[5\] net251 net726 vssd1 vssd1 vccd1 vccd1 _04739_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10700_ clknet_leaf_102_clk _00212_ net1162 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[172\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06686__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ clknet_leaf_32_clk _01192_ net1207 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06686__B2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08607__A _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06150__A3 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05894__C1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ clknet_leaf_93_clk _00143_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10562_ clknet_leaf_77_clk _00074_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10493_ net1497 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09388__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08060__B1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05949__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ clknet_leaf_111_clk _00626_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[586\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11045_ clknet_leaf_101_clk _00557_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[517\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06797__A _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10626__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07392__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05905__S net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__C net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09312__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06126__B1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11264__RESET_B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11878_ clknet_leaf_71_clk _01347_ net1271 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09112__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06772__S1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10829_ clknet_leaf_98_clk _00341_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09615__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07626__A0 _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09091__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05637__C1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06020_ core.register_file.registers_state\[875\] core.register_file.registers_state\[843\]
+ net667 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
XANTENNA__09379__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11401__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09067__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07971_ _03027_ _03402_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09710_ net243 net2474 net279 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
X_06922_ _03025_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08398__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07157__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__A0 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07155__X _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ net2352 net393 _05079_ net1002 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06853_ core.register_file.registers_state\[1007\] core.register_file.registers_state\[975\]
+ net853 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__mux2_1
XANTENNA__06500__A _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05804_ _01905_ _01906_ _01908_ _01907_ net648 net623 vssd1 vssd1 vccd1 vccd1 _01909_
+ sky130_fd_sc_hd__mux4_1
X_09572_ _04909_ net399 net301 net1965 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06784_ net1084 _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09303__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ core.pc.current_pc\[26\] core.pc.current_pc\[27\] _04583_ vssd1 vssd1 vccd1
+ vccd1 _04603_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05735_ net956 core.register_file.registers_state\[756\] net766 vssd1 vssd1 vccd1
+ vccd1 _01840_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout257_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06668__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ core.pc.current_pc\[20\] core.pc.current_pc\[21\] _04520_ vssd1 vssd1 vccd1
+ vccd1 _04540_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06668__B2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05666_ net1057 core.register_file.registers_state\[342\] vssd1 vssd1 vccd1 vccd1
+ _01771_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07405_ _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07331__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08385_ core.pc.current_pc\[14\] _04460_ net229 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05597_ net1042 core.register_file.registers_state\[219\] vssd1 vssd1 vccd1 vccd1
+ _01702_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout424_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1166_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire409 net410 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_128_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07336_ net1082 _03440_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08861__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09082__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07093__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__B _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ net1089 _03370_ _03371_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09006_ _04659_ _04758_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__nor2_1
XANTENNA__06840__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06218_ net625 _02321_ _02322_ _02320_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07198_ net1089 _03295_ _03296_ net967 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout793_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11081__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06149_ net947 core.register_file.registers_state\[455\] vssd1 vssd1 vccd1 vccd1
+ _02254_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__S net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06053__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net523 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_2
Xfanout531 net534 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_4
X_09908_ _05017_ net384 net375 net1661 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__a22o_1
Xfanout564 net566 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_2
Xfanout575 _04336_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_2
XANTENNA__09542__A0 _04887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07506__A _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_4
Xfanout597 net599 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_2
X_09839_ _04893_ net2153 net379 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10152__A1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06356__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11801_ clknet_leaf_54_clk _01302_ net1299 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08648__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11732_ clknet_leaf_45_clk _01244_ net1288 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07512__Y _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06409__X _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05867__C1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11663_ clknet_leaf_45_clk _01175_ net1288 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10614_ clknet_leaf_44_clk _00126_ net1286 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05882__A2 _01978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ clknet_leaf_27_clk _01106_ net1203 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05619__C1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10545_ clknet_leaf_76_clk _00057_ net1260 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10657__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08072__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10476_ net1370 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09781__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08800__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902__1319 vssd1 vssd1 vccd1 vccd1 _11902__1319/HI net1319 sky130_fd_sc_hd__conb_1
X_11028_ clknet_leaf_51_clk _00540_ net1297 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[500\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10143__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__X _03808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06362__A3 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05520_ _01490_ _01623_ _01624_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05858__C1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05451_ net1043 core.register_file.registers_state\[989\] core.register_file.registers_state\[1021\]
+ net672 net1011 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08170_ net1113 _04272_ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__o21ai_1
X_05382_ net967 _01483_ _01486_ net768 _01480_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__a311o_2
XFILLER_0_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07121_ net989 core.register_file.registers_state\[325\] net876 core.register_file.registers_state\[357\]
+ net1075 vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06822__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07052_ net990 core.register_file.registers_state\[455\] net876 core.register_file.registers_state\[487\]
+ net982 vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__a221o_1
XANTENNA__06822__B2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06003_ net1049 core.register_file.registers_state\[460\] vssd1 vssd1 vccd1 vccd1
+ _02108_ sky130_fd_sc_hd__or2_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XANTENNA__10017__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09772__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput189 net189 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__10941__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07954_ _04056_ _04058_ net485 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09524__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ _03004_ _03009_ net780 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07885_ net513 _03854_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout374_A _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ net743 _04995_ net459 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__and3_1
XANTENNA__06889__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06836_ net1087 _02939_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _04891_ net2145 net305 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__mux2_1
X_06767_ _02866_ _02871_ net781 vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__mux2_1
XANTENNA__11115__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ _02535_ _04586_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__or2_1
XANTENNA__07838__B1 _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05718_ net719 _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06376__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ _05003_ net322 net264 net1954 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__a22o_1
X_06698_ net790 _02799_ _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_82_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08437_ _01868_ _04523_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05649_ net949 core.register_file.registers_state\[758\] net763 vssd1 vssd1 vccd1
+ vccd1 _01754_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout1071_X net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1169_X net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07996__A _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08368_ _04460_ _04461_ net229 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__or3b_1
XANTENNA__09055__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07319_ net1095 core.register_file.registers_state\[347\] core.register_file.registers_state\[379\]
+ net837 net979 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_22_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07066__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09259__Y _05046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08299_ _04396_ _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08802__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08163__Y _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11597__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ _05115_ net1565 net238 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ net1315 net1989 _01442_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__o21a_1
XANTENNA__08566__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ net120 net920 net909 net1545 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1304 net1305 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__clkbuf_4
Xfanout1315 net34 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__buf_2
XANTENNA__10361__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 _05025_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_4
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07236__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 _04883_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_4
XANTENNA__06329__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06140__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout383 net386 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout394 _05066_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09294__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ clknet_leaf_53_clk net1744 net1302 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05978__X _02083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ clknet_leaf_70_clk _01158_ net1275 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07057__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_1
XFILLER_0_123_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput36 gpio_in[10] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_11577_ clknet_leaf_29_clk _01089_ net1200 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[25\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_103_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput47 gpio_in[20] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 gpio_in[30] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06265__C1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05607__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10528_ clknet_leaf_53_clk _00040_ net1300 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold809 core.register_file.registers_state\[253\] vssd1 vssd1 vccd1 vccd1 net2128
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10964__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06280__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10459_ net1327 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08557__A1 _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09754__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09626__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06568__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10116__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05791__A1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ net452 _02873_ net444 net509 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__a31o_1
XANTENNA__07532__A2 _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ net825 _02724_ _02725_ net786 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09340_ _04978_ net418 net413 net1645 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a22o_1
X_06552_ net975 _02655_ _02656_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__or3_1
X_05503_ net1058 core.register_file.registers_state\[732\] core.register_file.registers_state\[764\]
+ net684 net1030 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ net2348 net222 net335 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06483_ net1036 core.register_file.registers_state\[216\] core.register_file.registers_state\[248\]
+ net670 net651 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__o221a_1
XANTENNA__06209__B _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08222_ _01623_ _01626_ _01624_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05434_ net1047 core.register_file.registers_state\[94\] core.register_file.registers_state\[126\]
+ net676 net640 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08705__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07048__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ _04096_ _04140_ _04215_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__and4_1
X_05365_ core.register_file.registers_state\[286\] core.register_file.registers_state\[318\]
+ core.register_file.registers_state\[414\] core.register_file.registers_state\[446\]
+ net876 net1075 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07104_ net974 _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__and2_1
XANTENNA__05400__Y _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _03387_ _03389_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__o21ai_1
X_05296_ _01391_ _01408_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__or2_4
XFILLER_0_31_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07035_ _03139_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1031_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08711__Y _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07608__X _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout491_A _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout589_A _05093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ net745 net613 net226 vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09970__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A2 _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _04029_ _04030_ _04039_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_127_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11574__Q core.decoder.inst\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05782__A1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05782__B2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ net510 _03689_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__nand2_1
XANTENNA__09512__A3 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09607_ net2521 net394 _05069_ net1000 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__a22o_1
X_06819_ net1093 core.register_file.registers_state\[173\] net833 core.register_file.registers_state\[141\]
+ net804 vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05534__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07799_ net488 _03903_ _03896_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout923_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1286_X net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ net223 net2083 net304 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10837__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ _04969_ net325 net263 net1943 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ clknet_leaf_103_clk _01012_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[972\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08615__A _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_93_clk_X clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11901__1318 vssd1 vssd1 vccd1 vccd1 _11901__1318/HI net1318 sky130_fd_sc_hd__conb_1
XFILLER_0_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ clknet_leaf_91_clk _00943_ net1246 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[903\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10356__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ clknet_leaf_79_clk _00874_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[834\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11749__Q net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ _05098_ net1536 net238 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06262__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ clknet_leaf_17_clk _00805_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[765\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09736__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ net1126 net1433 net911 _05230_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input52_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09200__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1103 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_4
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ net1697 net916 net906 core.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 _01211_
+ sky130_fd_sc_hd__a22o_1
Xfanout1123 core.control_logic.instruction\[4\] vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1134 net1179 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_2
XANTENNA__07762__A2 _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1145 net1146 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__clkbuf_2
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_2
Xfanout1167 net1179 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05773__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1179 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05773__B2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_clk_X clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06722__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08475__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10672__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10282__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09120__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11629_ clknet_leaf_49_clk _01141_ net1309 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10266__S _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06316__Y _02421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10034__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__X _04860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold606 core.register_file.registers_state\[553\] vssd1 vssd1 vccd1 vccd1 net1925
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 core.register_file.registers_state\[646\] vssd1 vssd1 vccd1 vccd1 net1936
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 core.register_file.registers_state\[811\] vssd1 vssd1 vccd1 vccd1 net1947
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 core.register_file.registers_state\[256\] vssd1 vssd1 vccd1 vccd1 net1958
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09727__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08840_ _04714_ _04882_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__or2_4
XANTENNA__09075__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08771_ net733 _04004_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__nor2_1
XANTENNA__11292__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05983_ _02086_ _02087_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__or2_1
XANTENNA__05764__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _01708_ _03446_ net548 _01665_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07653_ _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06604_ _02707_ _02708_ net794 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07584_ _02519_ _03660_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__nor2_2
XFILLER_0_125_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09323_ _04951_ net416 net331 net1788 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a22o_1
X_06535_ net790 _02636_ _02639_ net776 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout337_A _05046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1079_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ net2539 net339 _05042_ _05043_ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06466_ net936 core.register_file.registers_state\[952\] net760 net1009 vssd1 vssd1
+ vccd1 vccd1 _02571_ sky130_fd_sc_hd__o31a_1
XANTENNA__06654__S net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08205_ _03774_ _03817_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05417_ net1007 net747 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__nand2_8
XFILLER_0_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09185_ _04975_ net357 net425 net1576 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__a22o_1
XANTENNA__10029__X _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout504_A _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06397_ core.register_file.registers_state\[1\] net704 net644 _02501_ vssd1 vssd1
+ vccd1 vccd1 _02502_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06229__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1246_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09965__S net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _03904_ _04130_ net533 vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__mux2_1
X_05348_ wb.curr_state\[0\] _01377_ core.WRITE_I net1125 net2537 vssd1 vssd1 vccd1
+ vccd1 _00009_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_116_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11569__Q core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08067_ _04157_ _04164_ _04171_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__or3_4
XFILLER_0_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05279_ core.control_logic.instruction\[6\] core.control_logic.instruction\[5\] net1123
+ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__and3b_1
XFILLER_0_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09718__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ net1101 core.register_file.registers_state\[456\] core.register_file.registers_state\[488\]
+ net845 net1074 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout873_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11635__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05755__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net565 _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_86_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07514__A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ clknet_leaf_97_clk _00443_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[403\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ clknet_leaf_88_clk _00374_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[334\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11015__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ clknet_leaf_16_clk _00305_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[265\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06468__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10016__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11165__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11414_ clknet_leaf_42_clk _00926_ net1283 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[886\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05691__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08632__X _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11345_ clknet_leaf_74_clk _00857_ net1255 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[817\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06866__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11289__RESET_B net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09709__A0 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07395__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05443__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ clknet_leaf_101_clk _00788_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[748\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09185__A1 _04975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ net74 net920 vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10158_ wb.curr_state\[0\] net910 _01452_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__o21a_1
XANTENNA__05746__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05746__B2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 core.register_file.registers_state\[26\] vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10089_ core.pc.current_pc\[15\] net591 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09115__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07499__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__A2 _04018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06171__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06320_ core.register_file.registers_state\[544\] core.register_file.registers_state\[512\]
+ net692 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08999__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05879__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06251_ net951 core.register_file.registers_state\[676\] net765 vssd1 vssd1 vccd1
+ vccd1 _02356_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06182_ net652 _02284_ _02286_ net620 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__o211a_1
XANTENNA__10009__B _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 core.register_file.registers_state\[824\] vssd1 vssd1 vccd1 vccd1 net1722
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11658__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold414 core.register_file.registers_state\[769\] vssd1 vssd1 vccd1 vccd1 net1733
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold425 _01227_ vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold436 core.register_file.registers_state\[676\] vssd1 vssd1 vccd1 vccd1 net1755
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08702__B net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold447 core.register_file.registers_state\[440\] vssd1 vssd1 vccd1 vccd1 net1766
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold458 core.register_file.registers_state\[552\] vssd1 vssd1 vccd1 vccd1 net1777
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06631__C1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09941_ core.decoder.inst\[30\] core.CPU_DAT_O\[30\] net893 vssd1 vssd1 vccd1 vccd1
+ _01094_ sky130_fd_sc_hd__mux2_1
Xhold469 core.register_file.registers_state\[378\] vssd1 vssd1 vccd1 vccd1 net1788
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout905 _05242_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout916 net917 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout927 net931 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_4
XANTENNA__10025__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ _04951_ net384 net266 net1792 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__a22o_1
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_2
XANTENNA__07726__A2 _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1103 core.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ _03862_ _04868_ net732 vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__mux2_1
XANTENNA__05737__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1114 core.register_file.registers_state\[165\] vssd1 vssd1 vccd1 vccd1 net2433
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout287_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1125 core.register_file.registers_state\[55\] vssd1 vssd1 vccd1 vccd1 net2444
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 core.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
X_11900__1317 vssd1 vssd1 vccd1 vccd1 _11900__1317/HI net1317 sky130_fd_sc_hd__conb_1
Xhold1147 core.register_file.registers_state\[125\] vssd1 vssd1 vccd1 vccd1 net2466
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net608 net216 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__and2_1
X_05966_ net936 core.register_file.registers_state\[941\] net760 net1009 vssd1 vssd1
+ vccd1 vccd1 _02071_ sky130_fd_sc_hd__o31a_1
Xhold1158 core.register_file.registers_state\[599\] vssd1 vssd1 vccd1 vccd1 net2477
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 core.register_file.registers_state\[128\] vssd1 vssd1 vccd1 vccd1 net2488
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _03696_ _03772_ _03809_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__a21o_2
XANTENNA__05406__X _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08687__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ net569 _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__and2_1
X_05897_ _02000_ _02001_ net618 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1196_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10594__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ _01391_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_66_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08864__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06162__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08439__B1 _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ net498 _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout621_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _04925_ net416 net331 net1940 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__a22o_1
XANTENNA__05789__A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06518_ core.register_file.registers_state\[541\] core.register_file.registers_state\[573\]
+ net868 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08165__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07111__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07498_ _03601_ _03602_ net1085 vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__o21a_1
XANTENNA__09651__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ net560 _04828_ _05034_ net341 net2110 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06449_ core.register_file.registers_state\[281\] core.register_file.registers_state\[313\]
+ core.register_file.registers_state\[409\] core.register_file.registers_state\[441\]
+ net714 net1023 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09939__A0 core.decoder.inst\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09695__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_X net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06870__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09168_ _04944_ net352 net343 net2228 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout990_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08119_ net484 _03716_ _03726_ net490 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ net2221 net365 net358 _04827_ vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07965__A2 _04018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ clknet_leaf_6_clk _00642_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[602\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold970 core.register_file.registers_state\[588\] vssd1 vssd1 vccd1 vccd1 net2289
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold981 core.register_file.registers_state\[754\] vssd1 vssd1 vccd1 vccd1 net2300
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 core.register_file.registers_state\[172\] vssd1 vssd1 vccd1 vccd1 net2311
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ clknet_leaf_93_clk _00573_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[533\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10012_ net1590 net541 net520 _05106_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__a22o_1
XANTENNA__06925__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
X_10914_ clknet_leaf_78_clk _00426_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[386\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06153__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11894_ clknet_leaf_53_clk _01363_ net1300 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10845_ clknet_leaf_20_clk _00357_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05900__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10776_ clknet_leaf_5_clk _00288_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[248\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07102__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09642__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10252__A3 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11328_ clknet_leaf_56_clk _00840_ net1294 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[800\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11259_ clknet_leaf_22_clk _00771_ net1184 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[731\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07169__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06042__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07264__S0 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05820_ net723 _01910_ _01918_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__05881__B _01958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05814__S1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06392__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06392__B2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05751_ net1064 core.register_file.registers_state\[468\] vssd1 vssd1 vccd1 vccd1
+ _01856_ sky130_fd_sc_hd__or2_1
XANTENNA__07016__S0 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_8
X_08470_ _04535_ _04554_ _04545_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06144__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05682_ net1056 core.register_file.registers_state\[725\] vssd1 vssd1 vccd1 vccd1
+ _01787_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07421_ net1091 core.register_file.registers_state\[88\] core.register_file.registers_state\[120\]
+ net834 net802 vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07892__A1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05352__C1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07352_ core.register_file.registers_state\[90\] core.register_file.registers_state\[122\]
+ net866 vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__mux2_1
XANTENNA__09094__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09633__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05402__A core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06303_ net1062 core.register_file.registers_state\[611\] net754 _02407_ vssd1 vssd1
+ vccd1 vccd1 _02408_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08841__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07283_ _03289_ _03292_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__or2_1
XANTENNA__11480__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ net564 _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_113_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06234_ core.register_file.registers_state\[869\] core.register_file.registers_state\[837\]
+ net682 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09397__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold200 net186 vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold211 core.IO_mod.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
X_06165_ net1029 _02268_ _02269_ net1006 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a31o_1
Xhold222 _01203_ vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 core.ADR_I\[7\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold244 net140 vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 core.IO_mod.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
X_06096_ _02198_ _02200_ net1028 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__o21a_1
XANTENNA__05958__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold266 net144 vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 _01230_ vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08151__C _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05958__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold288 core.register_file.registers_state\[826\] vssd1 vssd1 vccd1 vccd1 net1607
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ net1114 core.CPU_DAT_O\[13\] net894 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
Xhold299 core.IO_mod.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net708 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout713 net715 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
Xfanout724 _01498_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_6
XANTENNA__08859__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1111_A core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net740 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1209_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout746 _04653_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_4
X_09855_ _04917_ net385 net266 net2009 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__a22o_1
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 net759 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
Xfanout768 net770 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__buf_4
XANTENNA_fanout571_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 net780 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_4
XANTENNA_fanout669_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net732 _04853_ _04854_ _04852_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_107_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06383__A1 core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06998_ net972 _03101_ _03102_ net1067 vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__o31a_1
X_09786_ _04748_ net385 net273 net1818 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06383__B2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10704__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11582__Q core.decoder.inst\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ net572 net608 _04795_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__and3_1
X_05949_ net1037 core.register_file.registers_state\[173\] net669 core.register_file.registers_state\[141\]
+ net637 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout836_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_64_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ net2271 net468 net438 _04738_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a22o_1
XANTENNA__06135__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09872__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10578__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ _03722_ _03723_ net507 vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__mux2_1
X_08599_ _04306_ _04673_ _04317_ _04004_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ clknet_leaf_106_clk _00142_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09085__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ clknet_leaf_84_clk _00073_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10234__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10492_ net1426 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05949__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11203__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ clknet_leaf_17_clk _00625_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[585\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11044_ clknet_leaf_80_clk _00556_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[516\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07020__C1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10170__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_X net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09312__A1 _04935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05921__S net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__A2 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07874__A1 _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09620__C net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ clknet_leaf_52_clk _01346_ net1304 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10828_ clknet_leaf_102_clk _00340_ net1162 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[300\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09615__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08823__A0 _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07626__A1 _03730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ clknet_leaf_91_clk _00271_ net1239 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[231\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06834__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09067__C net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06062__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07970_ net530 _04066_ _04073_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__a21o_1
X_06921_ _03023_ _03024_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__nor2_1
XANTENNA__05892__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06852_ core.register_file.registers_state\[879\] core.register_file.registers_state\[847\]
+ net853 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__mux2_1
X_09640_ net745 _05015_ net461 vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and3_1
XANTENNA__10303__A _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06365__B2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05803_ core.register_file.registers_state\[978\] core.register_file.registers_state\[1010\]
+ net706 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__mux2_1
X_09571_ _04907_ net402 net300 net1932 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__a22o_1
X_06783_ core.register_file.registers_state\[784\] core.register_file.registers_state\[816\]
+ core.register_file.registers_state\[912\] core.register_file.registers_state\[944\]
+ net869 net1073 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_102_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_47_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_102_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08522_ _04594_ _04602_ core.pc.current_pc\[26\] net595 vssd1 vssd1 vccd1 vccd1 _00034_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05734_ net1063 core.register_file.registers_state\[596\] core.register_file.registers_state\[628\]
+ net691 net648 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__o221a_1
XANTENNA__09854__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ core.pc.current_pc\[20\] net596 _04537_ _04539_ vssd1 vssd1 vccd1 vccd1 _00028_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05665_ core.register_file.registers_state\[278\] core.register_file.registers_state\[310\]
+ core.register_file.registers_state\[406\] core.register_file.registers_state\[438\]
+ net706 net1022 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07404_ _03506_ _03508_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__or2_1
XANTENNA__05403__Y _01508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08384_ core.pc.current_pc\[14\] _04460_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05596_ net1042 core.register_file.registers_state\[91\] vssd1 vssd1 vccd1 vccd1
+ _01701_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07335_ core.register_file.registers_state\[795\] core.register_file.registers_state\[827\]
+ core.register_file.registers_state\[923\] core.register_file.registers_state\[955\]
+ net867 net1071 vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10216__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08714__Y _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1061_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_A net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05628__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ net996 core.register_file.registers_state\[448\] net890 core.register_file.registers_state\[480\]
+ net984 vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__a221o_1
XANTENNA__06662__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ net2165 net429 _04976_ net436 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__a22o_1
XANTENNA__11226__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06217_ net944 core.register_file.registers_state\[197\] net703 core.register_file.registers_state\[229\]
+ net643 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07197_ net1089 _03297_ _03298_ _03301_ net1067 vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__a311o_1
XANTENNA__09909__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout205_X net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06148_ net950 core.register_file.registers_state\[327\] net1017 vssd1 vssd1 vccd1
+ vccd1 _02253_ sky130_fd_sc_hd__a21o_1
XANTENNA__11577__Q core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08730__X _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout786_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07250__C1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06079_ net1051 core.register_file.registers_state\[585\] core.register_file.registers_state\[617\]
+ net677 net925 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1114_X net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout510 net512 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11376__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
Xfanout532 net534 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
X_09907_ net1120 _05079_ net377 net1813 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__a22o_1
Xfanout543 _05096_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_2
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_4
XANTENNA_fanout953_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 net566 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_4
Xfanout576 _04336_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07002__C1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07506__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout587 _01505_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_4
X_09838_ net211 net1800 net381 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06356__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__B _02488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ net603 net205 net287 net257 net1622 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_38_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11800_ clknet_leaf_76_clk _01301_ net1260 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06108__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08177__X _04282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ clknet_leaf_45_clk _01243_ net1288 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10359__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11662_ clknet_leaf_45_clk _01174_ net1288 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09058__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06138__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ clknet_leaf_60_clk _00125_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05882__A3 _01985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ clknet_leaf_24_clk _01105_ net1185 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10544_ clknet_leaf_108_clk _00056_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06425__X _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06292__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ net1420 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09230__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07241__C1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08800__B _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10743__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ clknet_leaf_12_clk _00539_ net1172 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08741__C1 _04799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05555__C1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09297__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08528__A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07432__A _02534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09123__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06319__Y _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05450_ net1043 core.register_file.registers_state\[861\] core.register_file.registers_state\[893\]
+ net672 net926 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05381_ net809 _01484_ _01485_ net1086 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07120_ core.register_file.registers_state\[293\] core.register_file.registers_state\[261\]
+ core.register_file.registers_state\[421\] core.register_file.registers_state\[389\]
+ net849 net1075 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07051_ net990 core.register_file.registers_state\[327\] net881 core.register_file.registers_state\[359\]
+ net1076 vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07480__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11399__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06002_ net941 core.register_file.registers_state\[492\] net761 vssd1 vssd1 vccd1
+ vccd1 _02107_ sky130_fd_sc_hd__or3_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09646__X _05081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XANTENNA__08024__A1 _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09221__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__B _01893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07953_ _03706_ _03710_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__nand2_1
XANTENNA__05794__C1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A1 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ _03005_ _03006_ _03007_ _03008_ net819 net790 vssd1 vssd1 vccd1 vccd1 _03009_
+ sky130_fd_sc_hd__mux4_1
X_07884_ _02782_ _03987_ _02752_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ net2270 net391 _05073_ net998 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__a22o_1
X_06835_ net991 core.register_file.registers_state\[463\] net877 core.register_file.registers_state\[495\]
+ net982 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout367_A _04898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ net214 net2408 net305 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__mux2_1
X_06766_ _02867_ _02868_ _02869_ _02870_ net792 net812 vssd1 vssd1 vccd1 vccd1 _02871_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06657__S net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05561__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ _02535_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__and2_1
X_05717_ _01813_ _01816_ _01821_ net625 net635 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a221o_1
XANTENNA__07838__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06697_ net785 _02800_ _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__or3_1
X_09485_ _05001_ net325 net263 net1930 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1276_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09968__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05849__B1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08436_ _01868_ _04523_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__nand2_1
X_05648_ net1056 core.register_file.registers_state\[598\] core.register_file.registers_state\[630\]
+ net684 net645 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__o221a_1
XANTENNA__06510__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11155__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06510__B2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08367_ core.pc.current_pc\[12\] _04440_ core.pc.current_pc\[13\] vssd1 vssd1 vccd1
+ vccd1 _04461_ sky130_fd_sc_hd__a21oi_1
X_05579_ net1040 core.register_file.registers_state\[731\] vssd1 vssd1 vccd1 vccd1
+ _01684_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1064_X net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08799__C1 _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07318_ core.register_file.registers_state\[283\] core.register_file.registers_state\[315\]
+ core.register_file.registers_state\[411\] core.register_file.registers_state\[443\]
+ net866 net1072 vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_134_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08298_ _04395_ _02274_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__and2b_1
XANTENNA__09460__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06274__B1 _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ _03351_ _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07471__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10260_ net1125 net2130 net910 _05238_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06026__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07223__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ net1743 net918 net908 core.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 _01227_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06577__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06577__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1305 net1313 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__buf_2
XANTENNA__07517__A _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 _05031_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09515__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout351 net353 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_4
Xfanout362 _05024_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout373 _04883_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_89_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout384 net386 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout395 net404 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_4
XANTENNA__07804__X _03909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08067__B _04164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11714_ clknet_leaf_50_clk net1504 net1308 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11645_ clknet_leaf_50_clk _01157_ net1307 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07398__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11541__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ clknet_leaf_27_clk _01088_ net1197 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09451__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 gpio_in[11] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
XFILLER_0_123_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput48 gpio_in[21] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06265__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput59 gpio_in[31] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_10527_ clknet_leaf_33_clk _00039_ net1205 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07462__C1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06315__B net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10458_ net1429 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09203__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08557__A2 _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11691__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10389_ net1332 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09626__B _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06568__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09118__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05791__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06620_ net993 core.register_file.registers_state\[661\] core.register_file.registers_state\[693\]
+ net881 net810 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a221o_1
XANTENNA__05543__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09809__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06551_ net1106 core.register_file.registers_state\[604\] core.register_file.registers_state\[636\]
+ net850 net810 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05502_ net950 core.register_file.registers_state\[700\] net707 core.register_file.registers_state\[668\]
+ net962 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10639__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09270_ net2468 _04889_ net335 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__mux2_1
XANTENNA__11529__SET_B net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06482_ net1035 core.register_file.registers_state\[88\] core.register_file.registers_state\[120\]
+ net665 net636 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08221_ _01490_ _01623_ _01627_ _03741_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05433_ _01535_ _01537_ net622 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08705__B _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ _04155_ _04172_ _04243_ _04256_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__nor4_1
XFILLER_0_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05364_ core.decoder.inst\[19\] _01397_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09442__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload54_A clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05410__A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ core.register_file.registers_state\[805\] core.register_file.registers_state\[773\]
+ core.register_file.registers_state\[933\] core.register_file.registers_state\[901\]
+ net849 net1075 vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08083_ _03387_ _03389_ net528 vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08796__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05295_ _01403_ net1123 core.control_logic.instruction\[5\] vssd1 vssd1 vccd1 vccd1
+ _01410_ sky130_fd_sc_hd__or3b_2
XANTENNA__09993__B2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07034_ net768 _03138_ _03126_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__o21a_2
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06008__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07205__C1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1024_A core.decoder.inst\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06559__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ net613 net227 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__and2_1
XANTENNA__05767__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__Q core.IO_mod.input_reg\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _03935_ _04040_ net533 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08867__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07867_ _03824_ _03971_ net495 vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__mux2_2
XANTENNA__11414__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__B1 _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout749_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08720__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09606_ net743 _04969_ net459 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06818_ core.register_file.registers_state\[13\] core.register_file.registers_state\[45\]
+ net865 vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07798_ _03790_ _03869_ net476 vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09537_ net224 net2425 net304 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06749_ core.register_file.registers_state\[17\] core.register_file.registers_state\[49\]
+ net885 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout916_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09698__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09681__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09468_ _04967_ net323 net263 net2074 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08419_ _04507_ _04508_ net229 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ net2189 net207 net408 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11430_ clknet_leaf_99_clk _00942_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09433__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06416__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05320__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__A1 core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ clknet_leaf_101_clk _00873_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[833\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10312_ _02272_ net1698 net236 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
XANTENNA__10900__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11292_ clknet_leaf_42_clk _00804_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[764\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08631__A core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10243_ net83 net914 vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07247__A _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ net132 net918 net908 net1523 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__a22o_1
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input45_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1113 net1114 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_4
Xfanout1124 core.pc.current_pc\[24\] vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_2
Xfanout1135 net1136 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_4
Xfanout1146 net1153 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_2
Xfanout1157 net1167 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__clkbuf_2
Xfanout1168 net1169 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_4
Xfanout1179 net1314 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08172__B1 _03909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09672__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05694__D1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11628_ clknet_leaf_72_clk _01140_ net1269 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10034__B2 _05117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11559_ clknet_leaf_25_clk _01071_ net1185 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06789__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 core.register_file.registers_state\[246\] vssd1 vssd1 vccd1 vccd1 net1926
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06789__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold618 core.register_file.registers_state\[742\] vssd1 vssd1 vccd1 vccd1 net1937
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10641__RESET_B net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06760__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold629 core.register_file.registers_state\[627\] vssd1 vssd1 vccd1 vccd1 net1948
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05997__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05461__B2 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05749__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08770_ core.IO_mod.input_reg\[21\] _04683_ net730 vssd1 vssd1 vccd1 vccd1 _04824_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05982_ net1044 core.register_file.registers_state\[972\] core.register_file.registers_state\[1004\]
+ net673 net1013 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07721_ _03660_ _03825_ _03824_ net493 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07652_ _03754_ _03756_ net484 vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06174__C1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06713__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06713__B2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06603_ net1105 core.register_file.registers_state\[214\] core.register_file.registers_state\[246\]
+ net851 net825 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07583_ net533 _03685_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__nand2_4
X_06534_ net785 _02637_ _02638_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09322_ _04949_ net422 net334 net2155 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07620__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06477__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10273__B2 core.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06465_ net637 _02566_ _02567_ _02568_ _02569_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09253_ core.register_file.registers_state\[317\] net475 net544 vssd1 vssd1 vccd1
+ vccd1 _05043_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout232_A _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08204_ _03798_ _03833_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__nor2_1
X_05416_ net932 net760 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__nor2_4
XANTENNA__05411__Y _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09184_ _04973_ net354 net424 net1889 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__a22o_1
X_06396_ net946 core.register_file.registers_state\[33\] net766 vssd1 vssd1 vccd1
+ vccd1 _02501_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08154__C _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ net513 _04134_ _04239_ _03694_ _02384_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a2111o_1
X_05347_ wb.curr_state\[0\] core.READ_I _01378_ net1125 wb.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _00008_ sky130_fd_sc_hd__a32o_1
XANTENNA__07426__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1141_A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1239_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08066_ _03771_ _03797_ _04167_ _04170_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05278_ core.control_logic.instruction\[3\] core.control_logic.instruction\[2\] core.control_logic.instruction\[0\]
+ core.control_logic.instruction\[1\] vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_102_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05452__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ net1101 core.register_file.registers_state\[328\] core.register_file.registers_state\[360\]
+ net845 net980 vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout699_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05452__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06242__Y _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1027_X net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09194__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10205__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11588__RESET_B net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _04860_ net601 vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__nor2_1
XANTENNA__10804__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ net531 _03686_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ net223 net737 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07514__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10930_ clknet_leaf_67_clk _00442_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[402\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06704__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05315__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ clknet_leaf_0_clk _00373_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[333\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10954__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09654__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10792_ clknet_leaf_14_clk _00304_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[264\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10367__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08209__A1 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07680__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05691__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09957__A1 core.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ clknet_leaf_63_clk _00925_ net1249 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07676__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11344_ clknet_leaf_104_clk _00856_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[816\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06866__S1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06640__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275_ clknet_leaf_107_clk _00787_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09185__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ net1127 net1474 net912 _05221_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07196__A1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10157_ net34 net1367 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__or2_1
XANTENNA__06943__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 core.register_file.registers_state\[956\] vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10088_ net472 _05151_ _05152_ net517 net1474 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09488__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10131__A _03964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06171__A2 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08448__A1 _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08095__X _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06250_ core.register_file.registers_state\[516\] net709 net646 _02354_ vssd1 vssd1
+ vccd1 vccd1 _02355_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09948__A1 core.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06181_ net1044 core.register_file.registers_state\[230\] net761 _02285_ net924 vssd1
+ vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_41_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold404 core.register_file.registers_state\[42\] vssd1 vssd1 vccd1 vccd1 net1723
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 core.register_file.registers_state\[301\] vssd1 vssd1 vccd1 vccd1 net1734
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold426 core.register_file.registers_state\[541\] vssd1 vssd1 vccd1 vccd1 net1745
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 core.register_file.registers_state\[805\] vssd1 vssd1 vccd1 vccd1 net1756
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05434__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold448 core.register_file.registers_state\[904\] vssd1 vssd1 vccd1 vccd1 net1767
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 core.ru.state\[3\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ core.decoder.inst\[29\] core.CPU_DAT_O\[29\] net894 vssd1 vssd1 vccd1 vccd1
+ _01093_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05434__B2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10827__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09176__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09871_ _04949_ net388 net268 net1993 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__a22o_1
Xfanout917 net921 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_2
Xfanout928 net931 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_2
XANTENNA__10025__B _01745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload17_A clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout939 net943 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_2
X_08822_ core.IO_mod.data_from_mem\[29\] core.IO_mod.input_reg\[29\] net250 vssd1
+ vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10191__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06395__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 core.register_file.registers_state\[95\] vssd1 vssd1 vccd1 vccd1 net2423
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06934__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1115 core.register_file.registers_state\[675\] vssd1 vssd1 vccd1 vccd1 net2434
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05834__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1126 core.register_file.registers_state\[166\] vssd1 vssd1 vccd1 vccd1 net2445
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 core.register_file.registers_state\[196\] vssd1 vssd1 vccd1 vccd1 net2456
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net733 _04298_ net526 _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__o211a_4
X_05965_ core.register_file.registers_state\[781\] core.register_file.registers_state\[813\]
+ net694 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
Xhold1148 core.register_file.registers_state\[315\] vssd1 vssd1 vccd1 vccd1 net2467
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 core.register_file.registers_state\[67\] vssd1 vssd1 vccd1 vccd1 net2478
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07704_ _03773_ _03788_ _03797_ _03808_ _03796_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a221o_1
X_05896_ net946 core.register_file.registers_state\[207\] net704 core.register_file.registers_state\[239\]
+ net644 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a221o_1
X_08684_ net605 _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09884__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ _01387_ _01492_ _01494_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__and3_2
XFILLER_0_95_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1091_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__Y _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1189_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__A1 _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07566_ net451 _03476_ net443 vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__and3_2
XANTENNA__10246__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ _04923_ net417 net332 net2232 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__a22o_1
XANTENNA__09100__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06517_ net973 _02620_ _02621_ net1066 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout235_X net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07111__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout614_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07497_ net1100 core.register_file.registers_state\[479\] core.register_file.registers_state\[511\]
+ net843 net1074 vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_118_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09236_ core.register_file.registers_state\[309\] net475 net545 vssd1 vssd1 vccd1
+ vccd1 _05034_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_79_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08880__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06448_ net648 _02547_ _02549_ net619 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06870__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09167_ _04942_ net358 net345 net1926 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__a22o_1
X_06379_ _01375_ _02475_ _02478_ _02483_ net634 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08118_ _03797_ _03922_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09098_ net2402 net365 net361 _04821_ vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout983_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05425__A1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ _03974_ _04017_ _04144_ _04149_ _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__o221a_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06413__B net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold960 core.register_file.registers_state\[695\] vssd1 vssd1 vccd1 vccd1 net2279
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 core.register_file.registers_state\[743\] vssd1 vssd1 vccd1 vccd1 net2290
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold982 core.register_file.registers_state\[704\] vssd1 vssd1 vccd1 vccd1 net2301
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ clknet_leaf_55_clk _00572_ net1295 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[532\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold993 core.register_file.registers_state\[712\] vssd1 vssd1 vccd1 vccd1 net2312
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _01502_ _01956_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__nor2_1
XANTENNA__10182__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07525__A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_103_clk_X clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913_ clknet_leaf_85_clk _00425_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[385\]
+ sky130_fd_sc_hd__dfrtp_1
X_11893_ clknet_leaf_72_clk _01362_ net1271 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11132__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10844_ clknet_leaf_40_clk _00356_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[316\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08356__A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07102__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10775_ clknet_leaf_22_clk _00287_ net1182 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06536__S0 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06310__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11282__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09618__C net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11327_ clknet_leaf_15_clk _00839_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[799\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05967__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09158__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11258_ clknet_leaf_6_clk _00770_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[730\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ net96 net920 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__and2_1
XANTENNA__07706__Y _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07264__S1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10173__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ clknet_leaf_94_clk _00701_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[661\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05507__X _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05750_ net956 core.register_file.registers_state\[500\] net765 vssd1 vssd1 vccd1
+ vccd1 _01855_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06129__C1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07016__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__X _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__X _03827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05681_ net1055 net753 core.register_file.registers_state\[789\] vssd1 vssd1 vccd1
+ vccd1 _01786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07420_ core.register_file.registers_state\[24\] core.register_file.registers_state\[56\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07892__A2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05352__B1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10228__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07351_ core.register_file.registers_state\[154\] core.register_file.registers_state\[186\]
+ net866 vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06302_ net954 core.register_file.registers_state\[579\] net1020 vssd1 vssd1 vccd1
+ vccd1 _02407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05402__B _01412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07282_ _03325_ _03385_ _03324_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06301__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06233_ core.register_file.registers_state\[805\] core.register_file.registers_state\[773\]
+ net682 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
X_09021_ net611 _04785_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06164_ net948 core.register_file.registers_state\[583\] net706 core.register_file.registers_state\[615\]
+ net659 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a221o_1
XANTENNA__09397__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 core.register_file.registers_state\[396\] vssd1 vssd1 vccd1 vccd1 net1520
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 net165 vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06514__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold223 core.register_file.registers_state\[414\] vssd1 vssd1 vccd1 vccd1 net1542
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08432__C _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06604__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold234 core.IO_mod.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06095_ net942 core.register_file.registers_state\[489\] net762 _02199_ net1015 vssd1
+ vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__o311a_1
Xhold245 core.register_file.registers_state\[33\] vssd1 vssd1 vccd1 vccd1 net1564
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 core.IO_mod.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 core.register_file.registers_state\[797\] vssd1 vssd1 vccd1 vccd1 net1586
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 net148 vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ core.decoder.inst\[12\] core.CPU_DAT_O\[12\] net892 vssd1 vssd1 vccd1 vccd1
+ _01076_ sky130_fd_sc_hd__mux2_1
XANTENNA__09149__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold289 net163 vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout703 net708 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_2
Xfanout714 net715 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__buf_4
XANTENNA__11109__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net731 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout397_A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 net740 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
Xfanout747 net752 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_8
X_09854_ _04915_ net386 net269 net1918 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__a22o_1
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06368__C1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1104_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_8
XANTENNA__07345__A _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ core.IO_mod.data_from_mem\[26\] net247 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_107_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _04743_ net390 net272 net1756 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ net1101 core.register_file.registers_state\[841\] core.register_file.registers_state\[873\]
+ net845 net980 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout564_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08736_ net610 net219 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__and2_1
X_05948_ net1112 net897 _01867_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a21o_1
XANTENNA__05591__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ net572 net608 net223 vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05879_ net634 _01974_ _01977_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout829_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10744__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ net449 net441 _03172_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09609__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ _04042_ _04278_ _04286_ _04298_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__or4b_1
XANTENNA__06540__C1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05894__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07549_ _03643_ _03653_ net480 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10560_ clknet_leaf_53_clk _00072_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06843__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _04748_ net417 net340 net1898 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10491_ net1373 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09388__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08060__A2 _03201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06071__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ clknet_leaf_13_clk _00624_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[584\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold790 core.register_file.registers_state\[439\] vssd1 vssd1 vccd1 vccd1 net2109
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11043_ clknet_leaf_66_clk _00555_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[515\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05582__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09312__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09863__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08086__A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ clknet_leaf_71_clk _01345_ net1274 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10827_ clknet_leaf_108_clk _00339_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10672__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07087__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08823__A1 _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ clknet_leaf_98_clk _00270_ net1160 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08814__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06834__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05637__B2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ clknet_leaf_84_clk _00201_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[161\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09379__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06062__A1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09645__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06920_ _03023_ _03024_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and2_1
XANTENNA__10146__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ core.register_file.registers_state\[815\] core.register_file.registers_state\[783\]
+ net853 vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__mux2_1
XANTENNA__10303__B _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05802_ core.register_file.registers_state\[850\] core.register_file.registers_state\[882\]
+ net712 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__mux2_1
X_09570_ _04905_ net401 net300 net2161 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__a22o_1
X_06782_ net771 _02881_ _02886_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_102_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08521_ net228 _04600_ _04601_ net595 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_102_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09303__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05733_ net662 _01836_ _01837_ net1032 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a31o_1
X_08452_ net208 _04538_ net596 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__o21ai_1
X_05664_ _01765_ _01766_ _01767_ _01768_ net625 net645 vssd1 vssd1 vccd1 vccd1 _01769_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06522__C1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07403_ _02561_ _03507_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08383_ _04472_ _04474_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__xnor2_1
X_05595_ net937 core.register_file.registers_state\[123\] net758 vssd1 vssd1 vccd1
+ vccd1 _01700_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07334_ net803 _03437_ _03438_ net1082 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08724__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07265_ net996 core.register_file.registers_state\[320\] net889 core.register_file.registers_state\[352\]
+ net1081 vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout312_A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09004_ net569 _04975_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06216_ net947 core.register_file.registers_state\[69\] net703 core.register_file.registers_state\[101\]
+ net657 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ net830 _03299_ _03300_ net976 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06244__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06147_ net1055 core.register_file.registers_state\[359\] net753 vssd1 vssd1 vccd1
+ vccd1 _02252_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_93_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07250__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06078_ net1051 core.register_file.registers_state\[713\] core.register_file.registers_state\[745\]
+ net678 net1015 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__o221a_1
XANTENNA__09790__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout500 net503 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_2
XANTENNA_fanout681_A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout779_A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout522 net524 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_2
X_09906_ _05014_ net384 net375 net2297 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__a22o_1
Xfanout533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_4
XFILLER_0_10_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1107_X net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_4
Xfanout555 _01506_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_8
Xfanout566 _04668_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_2
Xfanout577 _04336_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
XANTENNA__10996__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ net212 net1998 net379 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__mux2_1
Xfanout588 _05093_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10213__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 net600 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout946_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05307__B net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10925__RESET_B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _05005_ net293 net258 net1649 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08719_ net568 net607 net206 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09699_ net215 net2461 net279 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XANTENNA__08618__B _04306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11730_ clknet_leaf_37_clk _01242_ net1288 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07522__B _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06419__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05867__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05867__B2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ clknet_leaf_37_clk _01173_ net1222 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09058__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ clknet_leaf_53_clk _00124_ net1302 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11592_ clknet_leaf_33_clk _01104_ net1204 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08193__X _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08634__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06816__B1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05619__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10543_ clknet_leaf_83_clk _00055_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06292__A1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11768__Q core.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ net1393 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07241__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__A2 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10128__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11026_ clknet_leaf_68_clk _00538_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[498\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08741__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06752__C1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09404__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07713__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09297__A1 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08528__B _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07432__B _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06504__C1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05858__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05858__B2 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11859_ clknet_leaf_28_clk net55 net1196 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05380_ net988 core.register_file.registers_state\[702\] net870 core.register_file.registers_state\[670\]
+ net819 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__o221a_1
XANTENNA__06763__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07050_ core.register_file.registers_state\[295\] core.register_file.registers_state\[263\]
+ core.register_file.registers_state\[423\] core.register_file.registers_state\[391\]
+ net849 net1076 vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__mux4_1
XANTENNA__05379__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06064__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06001_ net1049 core.register_file.registers_state\[332\] core.register_file.registers_state\[364\]
+ net675 net925 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XANTENNA__08024__A2 _04018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__09221__A1 _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XANTENNA__09772__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07952_ _03706_ _03710_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__and2_1
XANTENNA__06991__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05408__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ core.register_file.registers_state\[972\] core.register_file.registers_state\[1004\]
+ net869 vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ _02752_ _02782_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__nand3_1
XFILLER_0_138_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06969__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ net742 _04993_ net457 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06834_ net991 core.register_file.registers_state\[335\] net877 core.register_file.registers_state\[367\]
+ net1077 vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a221o_1
XANTENNA__08719__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ net215 net2464 net306 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__mux2_1
XANTENNA__09288__A1 _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06765_ core.register_file.registers_state\[849\] core.register_file.registers_state\[881\]
+ net886 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A _05059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ core.pc.current_pc\[25\] _03506_ net574 vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__mux2_1
X_05716_ net645 _01817_ _01818_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a31o_1
X_09484_ _04999_ net318 net261 net1974 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__a22o_1
XANTENNA__06239__A core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ net1097 core.register_file.registers_state\[211\] core.register_file.registers_state\[243\]
+ net840 net819 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07394__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08435_ _01382_ net550 net575 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05647_ net928 _01750_ _01751_ net962 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ core.pc.current_pc\[12\] core.pc.current_pc\[13\] _04440_ vssd1 vssd1 vccd1
+ vccd1 _04460_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05578_ net1040 core.register_file.registers_state\[603\] vssd1 vssd1 vccd1 vccd1
+ _01683_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08799__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07317_ _03417_ _03420_ _02690_ _03415_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08297_ _04396_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11195__RESET_B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1057_X net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06274__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10070__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ net477 _03321_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout896_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10358__A0 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07179_ core.register_file.registers_state\[931\] core.register_file.registers_state\[899\]
+ net855 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1224_X net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07223__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ net1503 net919 net909 core.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 _01226_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09763__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08620__C _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1306 net1312 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout330 _05055_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
Xfanout341 _05031_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_8
XANTENNA__05318__A _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_4
XANTENNA__09515__A2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 net366 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_8
Xfanout374 _04883_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_4
Xfanout385 net386 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06140__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout396 net404 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_4
XFILLER_0_9_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09279__A1 _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06149__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11713_ clknet_leaf_50_clk net1456 net1307 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08239__C1 _02488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11644_ clknet_leaf_50_clk _01156_ net1307 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11575_ clknet_leaf_27_clk _01087_ net1197 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
XFILLER_0_108_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput38 gpio_in[12] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06265__A1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput49 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10526_ clknet_leaf_33_clk _00038_ net1205 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07462__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08651__X _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05473__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10349__A0 _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10457_ net1417 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09754__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09626__C net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ net1462 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05776__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06973__C1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10860__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ clknet_leaf_86_clk _00521_ net1226 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07714__Y _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05528__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06758__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06725__C1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08190__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05515__X _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05662__S net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06550_ net1104 core.register_file.registers_state\[732\] core.register_file.registers_state\[764\]
+ net850 net825 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05501_ net962 _01604_ _01605_ net659 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06481_ _02583_ _02585_ net620 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ _01625_ _04324_ _03742_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11366__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05432_ core.register_file.registers_state\[30\] net674 net654 _01536_ vssd1 vssd1
+ vccd1 vccd1 _01537_ sky130_fd_sc_hd__a211o_1
XANTENNA__06346__X _02451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05700__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08151_ _04186_ _04200_ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__nand3_1
X_05363_ core.decoder.inst\[19\] _01397_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__and2_4
XFILLER_0_28_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07102_ net989 core.register_file.registers_state\[837\] net875 core.register_file.registers_state\[869\]
+ net1075 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__a221o_1
XANTENNA__05410__B net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ _03826_ _04049_ net532 vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__mux2_1
X_05294_ net1123 core.control_logic.instruction\[5\] _01402_ vssd1 vssd1 vccd1 vccd1
+ _01409_ sky130_fd_sc_hd__and3b_4
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07033_ net968 _03132_ _03134_ _03137_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07618__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05409__Y _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08984_ _04704_ net2488 net429 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1017_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ _03983_ _04002_ _04013_ _04011_ net479 net495 vssd1 vssd1 vccd1 vccd1 _04040_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__05862__S0 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__A1 _01550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout477_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07866_ net476 _03925_ _03970_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06716__C1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08181__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ net2519 net394 _05068_ net1000 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__a22o_1
X_06817_ net970 _02918_ net775 vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07797_ core.decoder.inst\[24\] net898 net548 _03899_ _03901_ vssd1 vssd1 vccd1 vccd1
+ _03902_ sky130_fd_sc_hd__a221o_2
XANTENNA_fanout644_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09536_ net225 net2353 net304 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06748_ net1088 _02849_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08883__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09130__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ _04965_ net325 net263 net1866 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__a22o_1
X_06679_ net551 _02781_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A _01460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_A _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_X net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08418_ _04492_ _04496_ _04505_ _04506_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_93_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09398_ _04652_ _04654_ net604 _04710_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__nor4_2
XFILLER_0_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ _02117_ _04442_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06247__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05320__B net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11360_ clknet_leaf_57_clk _00872_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08912__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10311_ _02314_ net1469 net236 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ clknet_leaf_23_clk _00803_ net1186 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[763\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07087__X _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09197__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10883__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ net1126 net1440 net911 _05229_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09736__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__A1 core.decoder.inst\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10940__RESET_B net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1103 core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_4
X_10173_ net131 net916 net906 net1476 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1114 core.decoder.inst\[13\] vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__buf_4
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07815__X _03920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1136 net1140 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input38_A gpio_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1150 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11239__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1158 net1160 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_4
Xfanout1169 net1172 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08172__B2 _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08646__X _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05930__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07358__S0 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07132__C1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10282__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05511__A _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ clknet_leaf_70_clk _01139_ net1275 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09424__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10034__A2 _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire550 _02810_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_4
XFILLER_0_13_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11558_ clknet_leaf_25_clk _01070_ net1185 vssd1 vssd1 vccd1 vccd1 core.control_logic.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold608 core.register_file.registers_state\[140\] vssd1 vssd1 vccd1 vccd1 net1927
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10509_ clknet_leaf_45_clk _00021_ net1289 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold619 core.register_file.registers_state\[490\] vssd1 vssd1 vccd1 vccd1 net1938
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11489_ clknet_leaf_85_clk _01001_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[961\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09188__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09129__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05981_ net1044 core.register_file.registers_state\[844\] core.register_file.registers_state\[876\]
+ net673 net924 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07720_ net489 net476 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09360__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ net506 _03723_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06174__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06602_ net1105 core.register_file.registers_state\[86\] core.register_file.registers_state\[118\]
+ net851 net810 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__o221a_1
X_07582_ net512 _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nor2_1
XANTENNA__09112__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09321_ net558 _04947_ _05051_ net331 net2510 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
X_06533_ net1102 core.register_file.registers_state\[220\] core.register_file.registers_state\[252\]
+ net844 net822 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06477__A1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07620__B _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ net566 net559 _04871_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__and3_1
X_06464_ net943 core.register_file.registers_state\[696\] net747 net1009 vssd1 vssd1
+ vccd1 vccd1 _02569_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08203_ _02816_ _02845_ _04288_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__nand3_1
X_05415_ core.register_file.registers_state\[542\] core.register_file.registers_state\[574\]
+ net697 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__mux2_1
XANTENNA__09415__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09183_ _04971_ net354 net424 net1653 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__a22o_1
X_06395_ net1054 core.register_file.registers_state\[129\] net681 core.register_file.registers_state\[161\]
+ net658 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10039__A _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout225_A _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06229__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ net494 _04236_ _04238_ net533 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__o211a_1
XANTENNA__06229__B2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05346_ _01450_ _01452_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__nand2_1
XANTENNA__08623__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ _04017_ _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10769__RESET_B net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05277_ core.control_logic.instruction\[3\] core.control_logic.instruction\[2\] core.control_logic.instruction\[0\]
+ core.control_logic.instruction\[1\] vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__and4b_2
XFILLER_0_109_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1134_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09179__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ core.register_file.registers_state\[264\] core.register_file.registers_state\[296\]
+ core.register_file.registers_state\[392\] core.register_file.registers_state\[424\]
+ net872 net1074 vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_73_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09718__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout594_A _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1301_A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06937__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ net2148 net367 _04951_ net432 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ _03689_ _04018_ _04019_ _04021_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08898_ net2410 net369 _04905_ net438 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__a22o_1
XANTENNA__09351__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07849_ net1112 _03952_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__or2_1
XANTENNA__10221__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06165__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__C1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10860_ clknet_leaf_101_clk _00372_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[332\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05912__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07370__X _03475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ _04812_ net402 net309 net1872 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08001__S1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ clknet_leaf_92_clk _00303_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[263\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07022__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09406__A1 _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07680__A3 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10016__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ clknet_leaf_57_clk _00924_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[884\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05428__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11343_ clknet_leaf_83_clk _00855_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[815\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06640__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ clknet_leaf_0_clk _00786_ net1134 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[746\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11776__Q core.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10225_ net73 net920 vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__and2_1
XANTENNA__07815__S1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06928__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10115__C net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__X _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net2130 net515 _05200_ _05203_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05600__C1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 core.register_file.registers_state\[942\] vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10087_ _04268_ net590 vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__nand2_1
XANTENNA__08145__A1 _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06156__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload3_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__RESET_B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09412__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10989_ clknet_leaf_4_clk _00501_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[461\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06459__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05667__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06180_ net940 core.register_file.registers_state\[198\] vssd1 vssd1 vccd1 vccd1
+ _02285_ sky130_fd_sc_hd__and2_1
XANTENNA__07959__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11404__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold405 core.register_file.registers_state\[905\] vssd1 vssd1 vccd1 vccd1 net1724
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 core.register_file.registers_state\[916\] vssd1 vssd1 vccd1 vccd1 net1735
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold427 core.register_file.registers_state\[291\] vssd1 vssd1 vccd1 vccd1 net1746
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold438 core.register_file.registers_state\[874\] vssd1 vssd1 vccd1 vccd1 net1757
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06631__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold449 core.register_file.registers_state\[430\] vssd1 vssd1 vccd1 vccd1 net1768
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06631__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09870_ net558 _04947_ net456 net266 net1825 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__a32o_1
XANTENNA__09176__A3 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout907 _05205_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_2
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
Xfanout929 net931 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_8
X_08821_ net1957 net467 net434 _04867_ vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__a22o_1
XANTENNA__09581__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06395__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 core.register_file.registers_state\[722\] vssd1 vssd1 vccd1 vccd1 net2424
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 core.register_file.registers_state\[162\] vssd1 vssd1 vccd1 vccd1 net2435
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ core.IO_mod.data_from_mem\[18\] net246 _04808_ vssd1 vssd1 vccd1 vccd1 _04809_
+ sky130_fd_sc_hd__a21o_2
Xhold1127 core.register_file.registers_state\[204\] vssd1 vssd1 vccd1 vccd1 net2446
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 core.register_file.registers_state\[108\] vssd1 vssd1 vccd1 vccd1 net2457
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05964_ core.register_file.registers_state\[653\] core.register_file.registers_state\[685\]
+ net694 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
Xhold1149 core.register_file.registers_state\[330\] vssd1 vssd1 vccd1 vccd1 net2468
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ net489 _03802_ _03807_ _03664_ _03804_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a221o_1
XANTENNA__05416__A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09333__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ net733 _04155_ _04717_ _04750_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__o211ai_4
XANTENNA__08687__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05895_ net946 core.register_file.registers_state\[79\] net704 core.register_file.registers_state\[111\]
+ net658 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a221o_1
X_07634_ net255 _03738_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_105_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06698__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07631__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ net451 _03446_ net443 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08439__A2 _04511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout342_A _05031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09636__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _04921_ net416 net331 net1639 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1084_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06516_ net1096 core.register_file.registers_state\[861\] core.register_file.registers_state\[893\]
+ net837 net978 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ net1100 core.register_file.registers_state\[351\] core.register_file.registers_state\[383\]
+ net843 net980 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05658__C1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09235_ net560 _04822_ _05033_ net342 core.register_file.registers_state\[308\] vssd1
+ vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__a32o_1
X_06447_ _02550_ _02551_ net624 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06870__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ _04940_ net362 net345 net2004 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__a22o_1
X_06378_ _02479_ _02480_ _02482_ _02481_ net646 net623 vssd1 vssd1 vccd1 vccd1 _02483_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_75_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08117_ _04217_ _04219_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05329_ net1129 core.BUSY_O vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09097_ net2072 net363 net354 _04816_ vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08256__A_N net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08048_ _03730_ _03798_ _04150_ net547 _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__o221a_1
Xhold950 core.register_file.registers_state\[719\] vssd1 vssd1 vccd1 vccd1 net2269
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 core.register_file.registers_state\[208\] vssd1 vssd1 vccd1 vccd1 net2280
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout976_A _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05830__C1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 core.register_file.registers_state\[205\] vssd1 vssd1 vccd1 vccd1 net2291
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold983 core.register_file.registers_state\[322\] vssd1 vssd1 vccd1 vccd1 net2302
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1304_X net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold994 core.register_file.registers_state\[103\] vssd1 vssd1 vccd1 vccd1 net2313
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09572__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ net1648 net541 net520 _05105_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__a22o_1
XANTENNA__06710__A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _01498_ _02174_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and2_2
XANTENNA__11738__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06925__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10921__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09324__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10912_ clknet_leaf_55_clk _00424_ net1295 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[384\]
+ sky130_fd_sc_hd__dfrtp_1
X_11892_ clknet_leaf_49_clk _01361_ net1311 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06856__S net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10843_ clknet_leaf_21_clk _00355_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[315\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09627__B2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07638__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__A1_N net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ clknet_leaf_58_clk _00286_ net1286 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[246\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06536__S1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11577__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06074__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11326_ clknet_leaf_93_clk _00838_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[798\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11257_ clknet_leaf_55_clk _00769_ net1295 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[729\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09563__A0 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ net1128 net1655 net913 _05212_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a31o_1
XANTENNA__09407__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11188_ clknet_leaf_56_clk _00700_ net1295 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[660\]
+ sky130_fd_sc_hd__dfrtp_1
X_10139_ _05187_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08118__A1 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11408__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06129__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05680_ net1055 net753 core.register_file.registers_state\[917\] vssd1 vssd1 vccd1
+ vccd1 _01785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09142__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05352__B2 _01395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07350_ core.register_file.registers_state\[218\] core.register_file.registers_state\[250\]
+ net866 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__mux2_1
XANTENNA__08834__X _04878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06301_ net951 core.register_file.registers_state\[643\] net709 core.register_file.registers_state\[675\]
+ net646 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07281_ _03325_ _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__nor2_1
XANTENNA__06301__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09020_ net999 net463 _04986_ net428 net1927 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06232_ core.register_file.registers_state\[997\] core.register_file.registers_state\[965\]
+ net682 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06163_ net945 core.register_file.registers_state\[711\] net704 core.register_file.registers_state\[743\]
+ net643 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a221o_1
Xhold202 net169 vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09397__A3 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold213 net170 vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06065__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 net196 vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 core.register_file.registers_state\[897\] vssd1 vssd1 vccd1 vccd1 net1554
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 net188 vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
X_06094_ net1052 core.register_file.registers_state\[457\] vssd1 vssd1 vccd1 vccd1
+ _02199_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold257 core.register_file.registers_state\[263\] vssd1 vssd1 vccd1 vccd1 net1576
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 core.CPU_DAT_I\[13\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10944__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09922_ core.decoder.inst\[11\] core.CPU_DAT_O\[11\] net892 vssd1 vssd1 vccd1 vccd1
+ _01075_ sky130_fd_sc_hd__mux2_1
Xhold279 net184 vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout704 net708 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09554__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
Xfanout726 net731 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout737 net740 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
X_09853_ _04913_ net388 net267 net2273 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__a22o_1
XANTENNA__10164__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06530__A _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06368__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_2
XANTENNA_fanout292_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ core.IO_mod.input_reg\[26\] net252 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__nand2_1
XANTENNA__05417__Y _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _04738_ net387 net271 net1790 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ net1101 core.register_file.registers_state\[969\] core.register_file.registers_state\[1001\]
+ net845 net1074 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_68_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09306__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ net728 _04793_ _04794_ _04792_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__o31a_4
XFILLER_0_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05947_ net585 _02051_ _02018_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_64_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1299_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08666_ net608 net223 vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__and2_1
X_05878_ _01979_ _01980_ _01982_ _01981_ net623 net660 vssd1 vssd1 vccd1 vccd1 _01983_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08457__A _02747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07361__A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07617_ _03201_ _03631_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__or2_1
XANTENNA__06766__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08597_ _03917_ _03944_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout724_A _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_X net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07548_ _03651_ _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09085__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08293__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07479_ net1087 _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ _04743_ net419 net340 net1677 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10490_ net1428 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09149_ _04906_ net359 net346 net2226 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09793__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08920__A net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11111_ clknet_leaf_65_clk _00623_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[583\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06071__A2 _02174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold780 core.register_file.registers_state\[483\] vssd1 vssd1 vccd1 vccd1 net2099
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09545__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold791 core.register_file.registers_state\[309\] vssd1 vssd1 vccd1 vccd1 net2110
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07095__X _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ clknet_leaf_78_clk _00554_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[514\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06359__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09848__A1 _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07859__B1 _03963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11875_ clknet_leaf_76_clk _01344_ net1261 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10826_ clknet_leaf_106_clk _00338_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[298\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10757_ clknet_leaf_92_clk _00269_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[229\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10091__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06834__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06295__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06615__A _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10688_ clknet_leaf_53_clk _00200_ net1300 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[160\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09629__C net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06047__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__A1 core.decoder.inst\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09784__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ clknet_leaf_2_clk _00821_ net1139 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07896__A1_N _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09536__A0 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09137__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06850_ _02951_ _02952_ _02954_ _02953_ net792 net812 vssd1 vssd1 vccd1 vccd1 _02955_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07733__X _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05801_ core.register_file.registers_state\[786\] core.register_file.registers_state\[818\]
+ net712 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06781_ net1084 _02882_ _02885_ net779 vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__o211a_1
X_08520_ _04588_ _04598_ _04599_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05732_ net955 core.register_file.registers_state\[692\] net765 vssd1 vssd1 vccd1
+ vccd1 _01837_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_102_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08451_ core.pc.current_pc\[20\] _04520_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__xnor2_1
X_05663_ core.register_file.registers_state\[86\] core.register_file.registers_state\[118\]
+ net707 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ net537 _02598_ _02534_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ _04455_ _04473_ _04472_ _04464_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__o211a_1
XANTENNA__11742__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05594_ _01697_ _01698_ net617 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09600__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ net987 core.register_file.registers_state\[699\] net867 core.register_file.registers_state\[667\]
+ net818 vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08724__B _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05628__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07264_ core.register_file.registers_state\[288\] core.register_file.registers_state\[256\]
+ core.register_file.registers_state\[416\] core.register_file.registers_state\[384\]
+ net858 net1081 vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09003_ _04659_ _04751_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nor2_2
X_06215_ _02317_ _02319_ net617 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07195_ net1111 core.register_file.registers_state\[674\] core.register_file.registers_state\[642\]
+ net856 net812 vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout305_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06146_ _02247_ _02250_ net629 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_93_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06589__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07250__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06077_ _02178_ _02181_ net933 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11122__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 net503 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout1214_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout512 _02422_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _05013_ net384 net375 net1544 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__a22o_1
Xfanout534 _02423_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
XFILLER_0_10_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout674_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _04708_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_8
Xfanout556 net557 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07002__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07002__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ net205 net2532 net379 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_4
Xfanout578 _03617_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout589 _05093_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06979_ _03080_ _03082_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11272__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _05003_ net293 net259 net1840 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout939_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08718_ net607 net206 vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__and2_1
X_09698_ net216 net2424 net280 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
XANTENNA__05604__A _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ core.IO_mod.data_from_mem\[2\] net249 _04721_ vssd1 vssd1 vccd1 vccd1 _04722_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10965__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07522__C _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06419__B _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ clknet_leaf_45_clk _01172_ net1288 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08915__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09058__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ clknet_leaf_97_clk _00123_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11591_ clknet_leaf_25_clk _01103_ net1186 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08634__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ clknet_leaf_82_clk _00054_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08018__B1 _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10473_ net1398 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06029__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09766__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09230__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__C1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07241__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09781__A3 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11615__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ clknet_leaf_73_clk _00537_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08741__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07553__X _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06201__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05555__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07713__B _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11765__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09297__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10635__RESET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11858_ clknet_leaf_29_clk net54 net1195 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08825__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09420__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10809_ clknet_leaf_68_clk _00321_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11789_ clknet_leaf_29_clk _01293_ net1200 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06268__C1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11485__SET_B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08009__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07480__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07480__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11145__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06000_ _02101_ _02104_ net632 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07728__X _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05491__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09757__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_71_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09509__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__inv_2
XANTENNA__06080__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05794__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11295__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05794__B2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06902_ core.register_file.registers_state\[844\] core.register_file.registers_state\[876\]
+ net869 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07882_ _02905_ _03412_ _02785_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__a21o_1
XANTENNA__05408__B net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_86_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ net2070 net394 _05072_ net1000 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__a22o_1
X_06833_ core.register_file.registers_state\[303\] core.register_file.registers_state\[271\]
+ core.register_file.registers_state\[431\] core.register_file.registers_state\[399\]
+ net847 net1076 vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux4_1
XANTENNA__06969__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08719__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ net216 net2400 net304 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__mux2_1
X_06764_ core.register_file.registers_state\[785\] core.register_file.registers_state\[817\]
+ net886 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__mux2_1
X_08503_ _04573_ _04578_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__or2_1
XANTENNA__07299__A1 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05715_ net949 core.register_file.registers_state\[245\] net753 _01819_ net1022 vssd1
+ vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__o2111a_1
X_09483_ _04997_ net324 net263 net1929 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__a22o_1
X_06695_ net1097 core.register_file.registers_state\[83\] core.register_file.registers_state\[115\]
+ net840 net805 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__o221a_1
XANTENNA__06239__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ _04520_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07394__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05646_ net1056 core.register_file.registers_state\[854\] vssd1 vssd1 vccd1 vccd1
+ _01751_ sky130_fd_sc_hd__or2_1
XANTENNA__06954__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ core.pc.current_pc\[12\] net597 _04457_ _04459_ vssd1 vssd1 vccd1 vccd1 _00020_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_138_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05577_ net937 core.register_file.registers_state\[635\] net758 vssd1 vssd1 vccd1
+ vccd1 _01682_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout422_A _05029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08799__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07316_ _02905_ _03412_ _03420_ _02786_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a211o_1
XANTENNA__06259__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08296_ core.decoder.inst\[27\] net734 _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10048__Y _05127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09460__A2 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07247_ _03351_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07471__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07471__B2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__Y _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ core.register_file.registers_state\[995\] core.register_file.registers_state\[963\]
+ net848 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout791_A _01455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07223__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06129_ net1047 core.register_file.registers_state\[168\] net678 core.register_file.registers_state\[136\]
+ net641 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a221o_1
XANTENNA__08420__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11164__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1307 net1312 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout320 net326 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout331 _05047_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_6
Xfanout342 _05031_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout353 net362 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_4
XANTENNA__09515__A3 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout364 net366 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_4
Xfanout375 net378 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09920__A0 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout386 _05085_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09819_ _04885_ net2146 net379 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout397 net404 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_4
XANTENNA__06734__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05605__Y _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08487__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11712_ clknet_leaf_49_clk net1489 net1309 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ clknet_leaf_49_clk _01155_ net1309 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05988__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09987__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ clknet_leaf_25_clk _01086_ net1191 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[22\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
X_10525_ clknet_leaf_33_clk _00037_ net1207 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput39 gpio_in[13] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07462__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09739__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ net1351 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09203__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07214__A1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ net1421 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__05776__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ clknet_leaf_51_clk _00520_ net1304 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09415__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05528__A1 core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10816__RESET_B net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05500_ net1058 core.register_file.registers_state\[604\] core.register_file.registers_state\[636\]
+ net683 net1030 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__o221a_1
XANTENNA__06489__C1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06480_ core.register_file.registers_state\[24\] net670 net652 _02584_ vssd1 vssd1
+ vccd1 vccd1 _02585_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05431_ net1047 core.register_file.registers_state\[62\] net750 vssd1 vssd1 vccd1
+ vccd1 _01536_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05250__Y _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ _04254_ _04247_ _04245_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__and3b_4
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05362_ net790 _01461_ net776 _01466_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09442__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07101_ net989 core.register_file.registers_state\[965\] net875 core.register_file.registers_state\[997\]
+ net982 vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__a221o_1
X_08081_ _03993_ _04017_ _04175_ _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__o211a_4
XFILLER_0_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05293_ _01364_ net1123 _01401_ _01404_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__o211a_4
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05464__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ net969 _03135_ _03136_ net1066 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__o31a_1
XANTENNA__06661__C1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07205__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07618__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10685__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05419__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06014__S net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05767__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ net1116 _04654_ net611 _04710_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__or4_1
XANTENNA__05767__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07934_ _03686_ _04038_ _04036_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__o21ai_2
XANTENNA__05862__S1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09902__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07865_ net476 _03968_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_88_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A _04883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ net743 _04967_ net459 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__and3_1
XANTENNA__06811__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06816_ _02919_ _02920_ net1083 vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__o21a_1
X_07796_ net1003 _03899_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_84_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09535_ net226 net2462 net305 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__mux2_1
X_06747_ net976 _02850_ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout637_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ _04963_ net321 net264 net1953 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__a22o_1
X_06678_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__inv_2
XANTENNA__07141__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08417_ _04492_ _04496_ _04505_ _04506_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__or4bb_1
X_05629_ _01731_ _01733_ net621 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a21o_1
X_09397_ net607 net241 net319 net328 net1636 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout804_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1167_X net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10028__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__inv_2
XANTENNA__08752__X _04809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09433__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06416__C net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ _04378_ _04379_ _04376_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08641__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05320__C core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _02343_ net1584 net238 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06652__C1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11290_ clknet_leaf_7_clk _00802_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[762\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ net82 net915 vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07747__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ net130 net917 net907 net1507 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1106 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_4
Xfanout1115 net1117 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_8
Xfanout1126 _01379_ vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_4
Xfanout1137 net1139 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1148 net1150 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_4
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08172__A2 _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07358__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05999__A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07132__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09672__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08880__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05694__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ clknet_leaf_72_clk _01138_ net1269 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11557_ clknet_leaf_25_clk _01069_ net1185 vssd1 vssd1 vccd1 vccd1 core.control_logic.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
Xwire551 _02778_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_4
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05446__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ clknet_leaf_45_clk _00020_ net1288 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold609 core.register_file.registers_state\[189\] vssd1 vssd1 vccd1 vccd1 net1928
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11488_ clknet_leaf_57_clk _01000_ net1296 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[960\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05997__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05997__B2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__RESET_B net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ net1385 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10145__A _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05749__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05749__B2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06946__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05980_ core.decoder.inst\[12\] net896 _01867_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a21o_2
XFILLER_0_40_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09360__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ net500 _03701_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06174__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08984__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06601_ core.register_file.registers_state\[22\] core.register_file.registers_state\[54\]
+ net880 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07581_ _02384_ _03684_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__or2_4
XFILLER_0_125_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09320_ core.register_file.registers_state\[376\] net474 net544 vssd1 vssd1 vccd1
+ vccd1 _05051_ sky130_fd_sc_hd__o21a_1
X_06532_ net1102 core.register_file.registers_state\[92\] core.register_file.registers_state\[124\]
+ net844 net806 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08285__A _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09663__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07123__B1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05702__A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ net2453 net340 _05041_ _04867_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__a22o_1
XANTENNA__08871__A0 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06463_ net1037 net752 core.register_file.registers_state\[664\] vssd1 vssd1 vccd1
+ vccd1 _02568_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_135_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07620__C net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08202_ _02845_ _04288_ _02816_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05414_ net941 core.register_file.registers_state\[670\] core.register_file.registers_state\[702\]
+ net698 net639 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09182_ _04969_ net359 net425 net1604 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__a22o_1
XANTENNA__06009__S net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06394_ _02491_ _02492_ _02496_ _02498_ net963 net934 vssd1 vssd1 vccd1 vccd1 _02499_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05780__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10039__B _01549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08133_ net484 _04211_ _04237_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05345_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__inv_2
XANTENNA__07426__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__B1 _04691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07426__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout218_A _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05437__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08064_ _03791_ _04168_ net531 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__mux2_1
XANTENNA__06634__C1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05276_ _01388_ _01390_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ net790 _03116_ _03119_ net776 vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1127_A _01379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout587_A _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08966_ net565 _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07917_ _02385_ _03694_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net572 net224 net737 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout754_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
X_07848_ net546 _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__nor2_1
XANTENNA__06165__A1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__X _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05912__A1 core.decoder.inst\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05373__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ net527 _03813_ _03863_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__o31a_2
XANTENNA__11826__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09518_ _04807_ net400 net309 net1893 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__a22o_1
X_10790_ clknet_leaf_101_clk _00302_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[262\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09654__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__A1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ _04932_ net323 net314 net2294 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10850__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08923__A _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05771__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11411_ clknet_leaf_10_clk _00923_ net1149 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[883\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05691__A3 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11342_ clknet_leaf_89_clk _00854_ net1235 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[814\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05979__A1 _02083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06443__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11273_ clknet_leaf_38_clk _00785_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[745\]
+ sky130_fd_sc_hd__dfrtp_1
X_10224_ net1127 net1602 net912 _05220_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__a31o_1
XANTENNA_input50_A gpio_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ net556 _05201_ _05202_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07028__S0 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10086_ core.pc.current_pc\[14\] net592 vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__or2_1
Xhold6 core.register_file.registers_state\[996\] vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08145__A2 _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06156__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10988_ clknet_leaf_101_clk _00500_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[460\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05522__A _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07213__S net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06459__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08853__A0 _04887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07751__S1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11609_ clknet_leaf_29_clk _01121_ net1200 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06616__C1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06353__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 core.register_file.registers_state\[812\] vssd1 vssd1 vccd1 vccd1 net1725
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 core.register_file.registers_state\[807\] vssd1 vssd1 vccd1 vccd1 net1736
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 core.register_file.registers_state\[523\] vssd1 vssd1 vccd1 vccd1 net1747
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold439 core.register_file.registers_state\[793\] vssd1 vssd1 vccd1 vccd1 net1758
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_4
Xfanout919 net921 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_2
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ net570 net610 net210 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06395__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10191__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 core.register_file.registers_state\[579\] vssd1 vssd1 vccd1 vccd1 net2425
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 core.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ core.IO_mod.input_reg\[18\] net250 net725 vssd1 vssd1 vccd1 vccd1 _04808_
+ sky130_fd_sc_hd__a21o_1
Xhold1128 core.register_file.registers_state\[66\] vssd1 vssd1 vccd1 vccd1 net2447
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05963_ core.register_file.registers_state\[525\] net694 net636 vssd1 vssd1 vccd1
+ vccd1 _02068_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_77_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10723__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1139 core.register_file.registers_state\[72\] vssd1 vssd1 vccd1 vccd1 net2458
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09333__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07702_ _03805_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__and2b_1
XANTENNA__05416__B net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08682_ core.IO_mod.data_from_mem\[7\] net247 _04749_ vssd1 vssd1 vccd1 vccd1 _04750_
+ sky130_fd_sc_hd__a21o_2
X_05894_ net644 _01996_ _01998_ net625 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_120_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09884__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07912__A _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07895__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07633_ _03735_ _03736_ _03737_ net537 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_105_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05355__C1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07564_ net493 _03666_ _03668_ net513 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__a31o_1
XANTENNA__07631__B net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09097__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06528__A _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09636__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06515_ net1096 core.register_file.registers_state\[989\] core.register_file.registers_state\[1021\]
+ net837 net1070 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__o221a_1
X_09303_ _04919_ net416 net331 net1966 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__a22o_1
XANTENNA__08844__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10246__A3 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07495_ core.register_file.registers_state\[287\] core.register_file.registers_state\[319\]
+ core.register_file.registers_state\[415\] core.register_file.registers_state\[447\]
+ net873 core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_A _05046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1077_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06446_ net1064 core.register_file.registers_state\[217\] core.register_file.registers_state\[249\]
+ net690 net663 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__o221a_1
X_09234_ core.register_file.registers_state\[308\] _04666_ net545 vssd1 vssd1 vccd1
+ vccd1 _05033_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06962__S net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08743__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11229__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09165_ _04938_ net360 net346 net2361 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__a22o_1
X_06377_ core.register_file.registers_state\[994\] core.register_file.registers_state\[962\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout502_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1244_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08116_ net1113 _04218_ _04220_ net579 vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__o211a_1
X_05328_ net1129 core.BUSY_O vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__nor2_1
X_09096_ net2238 net365 net360 _04811_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06083__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08047_ net1112 _04150_ _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05259_ net1055 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XANTENNA__10919__RESET_B net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold940 core.register_file.registers_state\[71\] vssd1 vssd1 vccd1 vccd1 net2259
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold951 core.register_file.registers_state\[656\] vssd1 vssd1 vccd1 vccd1 net2270
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold962 core.register_file.registers_state\[581\] vssd1 vssd1 vccd1 vccd1 net2281
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 core.register_file.registers_state\[249\] vssd1 vssd1 vccd1 vccd1 net2292
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 core.register_file.registers_state\[501\] vssd1 vssd1 vccd1 vccd1 net2303
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 core.register_file.registers_state\[193\] vssd1 vssd1 vccd1 vccd1 net2314
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09998_ net1523 net542 net521 _05099_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__a22o_1
XANTENNA__10182__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ net2471 net370 _04939_ net439 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09875__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ clknet_leaf_16_clk _00423_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[383\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11891_ clknet_leaf_50_clk _01360_ net1307 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__A2_N _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05897__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__B _02717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09088__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ clknet_leaf_9_clk _00354_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[314\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05992__S0 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09627__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05342__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10773_ clknet_leaf_60_clk _00285_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[245\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11360__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08653__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06310__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05488__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07269__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11787__Q core.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07810__A1 _03697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07271__C1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11325_ clknet_leaf_19_clk _00837_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[797\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ clknet_leaf_4_clk _00768_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[728\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07023__C1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ net95 net919 vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__and2_1
X_11187_ clknet_leaf_98_clk _00699_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[659\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10173__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ core.pc.current_pc\[29\] _05183_ _05092_ vssd1 vssd1 vccd1 vccd1 _05188_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__05517__A core.decoder.inst\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10069_ _04155_ net557 net591 core.pc.current_pc\[7\] net472 vssd1 vssd1 vccd1 vccd1
+ _05141_ sky130_fd_sc_hd__o221a_1
XANTENNA__06129__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__B1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07877__A1 _03650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07877__B2 _03730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05888__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09079__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10228__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06300_ core.register_file.registers_state\[515\] net687 net660 _02404_ vssd1 vssd1
+ vccd1 vccd1 _02405_ sky130_fd_sc_hd__a211o_1
X_07280_ _03383_ _03384_ _03354_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06301__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11030__RESET_B net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06231_ core.register_file.registers_state\[933\] core.register_file.registers_state\[901\]
+ net682 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08054__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06162_ net658 _02265_ _02266_ net963 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_clk_X clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 core.register_file.registers_state\[801\] vssd1 vssd1 vccd1 vccd1 net1522
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 core.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06093_ net942 core.register_file.registers_state\[361\] net762 _02197_ net925 vssd1
+ vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__o311a_1
Xhold225 core.register_file.registers_state\[922\] vssd1 vssd1 vccd1 vccd1 net1544
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 core.register_file.registers_state\[781\] vssd1 vssd1 vccd1 vccd1 net1555
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold247 net149 vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold258 core.register_file.registers_state\[43\] vssd1 vssd1 vccd1 vccd1 net1577
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net1116 core.CPU_DAT_O\[10\] net892 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__mux2_1
Xhold269 _01214_ vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout705 net708 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11671__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 _01513_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_4
Xfanout727 net731 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
X_09852_ _04911_ net385 net269 net1883 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__a22o_1
Xfanout738 net740 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06368__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 net752 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_4
X_08803_ net727 _03884_ net525 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__a21o_1
XANTENNA__05576__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09783_ _04732_ net389 net271 net1694 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__a22o_1
X_06995_ net1085 _03099_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout285_A _05081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07913__Y _04018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ core.IO_mod.data_from_mem\[15\] net246 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__and2_2
XANTENNA__06957__S net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05946_ _02035_ _02036_ _02044_ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__o22ai_4
XANTENNA__05591__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _04734_ _04735_ _04733_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a21oi_4
X_05877_ core.register_file.registers_state\[913\] core.register_file.registers_state\[945\]
+ net711 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__mux2_1
XANTENNA__07412__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07616_ _03717_ _03720_ net483 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08596_ _03916_ _03943_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__nor2_1
XANTENNA__06540__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09609__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11051__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ net502 _03645_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout717_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10619__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08293__A1 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ core.register_file.registers_state\[799\] core.register_file.registers_state\[831\]
+ core.register_file.registers_state\[927\] core.register_file.registers_state\[959\]
+ net873 net1077 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__mux4_1
XANTENNA__09490__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09217_ _04738_ net421 net341 net1763 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06429_ _02532_ _02533_ _01632_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05500__C1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09148_ _04904_ net360 net346 net2342 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__B net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07253__C1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ net2218 net365 net357 _04720_ vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__a22o_1
XANTENNA__06151__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08920__B net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ clknet_leaf_98_clk _00622_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[582\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 core.register_file.registers_state\[485\] vssd1 vssd1 vccd1 vccd1 net2089
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold781 core.register_file.registers_state\[869\] vssd1 vssd1 vccd1 vccd1 net2100
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ clknet_leaf_85_clk _00553_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[513\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold792 core.register_file.registers_state\[259\] vssd1 vssd1 vccd1 vccd1 net2111
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__B net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__C1 _04809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06867__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07552__A _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11874_ clknet_leaf_72_clk _01343_ net1271 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10825_ clknet_leaf_40_clk _00337_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[297\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06819__C1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08284__A1 _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ clknet_leaf_77_clk _00268_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06455__X _02560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10091__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07492__C1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ clknet_leaf_14_clk _00199_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[159\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09233__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09784__A1 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09418__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ clknet_leaf_103_clk _00820_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[780\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08322__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11239_ clknet_leaf_65_clk _00751_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[711\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07446__B net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05800_ core.register_file.registers_state\[914\] core.register_file.registers_state\[946\]
+ net712 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__mux2_1
X_06780_ net971 _02883_ _02884_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05731_ net1063 net755 core.register_file.registers_state\[660\] vssd1 vssd1 vccd1
+ vccd1 _01836_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_102_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11074__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05253__Y _01368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08450_ net228 _04535_ _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__nor3_1
X_05662_ core.register_file.registers_state\[22\] core.register_file.registers_state\[54\]
+ net706 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06522__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05956__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06522__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11211__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07401_ _03494_ _03505_ net774 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__mux2_8
X_08381_ _04455_ _04473_ _04464_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__o21ai_1
X_05593_ net938 core.register_file.registers_state\[155\] net758 net922 vssd1 vssd1
+ vccd1 vccd1 _01698_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07332_ core.register_file.registers_state\[539\] core.register_file.registers_state\[571\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__mux2_1
XANTENNA__08275__A1 _03231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09472__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07401__S net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06286__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07263_ _01372_ _03360_ _03367_ net769 vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__a211oi_2
XANTENNA__10911__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07483__C1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09002_ net2306 net428 _04974_ net433 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__a22o_1
X_06214_ core.register_file.registers_state\[5\] net698 net639 _02318_ vssd1 vssd1
+ vccd1 vccd1 _02319_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07194_ core.register_file.registers_state\[546\] core.register_file.registers_state\[514\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__mux2_1
XANTENNA__09224__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__X _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06145_ net625 _02248_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__and3_1
XANTENNA__09775__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07786__A0 _03889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06076_ net960 _02179_ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__or3_1
XANTENNA__06541__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_2
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09904_ net1120 _05011_ net460 net377 net1547 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__a32o_1
Xfanout513 _02422_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1207_A net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
Xfanout557 _05091_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_4
X_09835_ net213 net1785 net380 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05549__C1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 _04668_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_4
Xfanout579 _03617_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout667_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _05001_ net297 net259 net1912 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06978_ _03080_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nand2_1
XANTENNA__05564__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07372__A _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05444__X _01549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ net525 _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__nor2_2
XFILLER_0_94_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05929_ net657 _02031_ _02032_ _02033_ net1006 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a311o_1
X_09697_ net217 net2174 net280 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout834_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08187__B _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08648_ core.IO_mod.input_reg\[2\] net253 net729 vssd1 vssd1 vccd1 vccd1 _04721_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08755__X _04812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07522__D _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06419__C _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08579_ net1121 net895 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10610_ clknet_leaf_70_clk _00122_ net1275 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11590_ clknet_leaf_27_clk _01102_ net1197 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05620__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10541_ clknet_leaf_98_clk _00053_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08018__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09215__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ net1357 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06029__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08650__B _04215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07529__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__X _03939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ clknet_leaf_105_clk _00536_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[496\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11097__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06201__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08741__A2 _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__A _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05354__X _01459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__B2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_X net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06504__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06504__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11857_ clknet_leaf_28_clk net53 net1195 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10808_ clknet_leaf_10_clk _00320_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09454__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11788_ clknet_leaf_28_clk _01292_ net1196 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06268__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10739_ clknet_leaf_12_clk _00251_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[211\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10148__A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06363__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08009__A1 _02206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09206__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA__06361__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__A1 _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ _03699_ _03709_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06991__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ core.register_file.registers_state\[908\] core.register_file.registers_state\[940\]
+ net869 vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
X_07881_ _02905_ _03412_ _02785_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08193__B1 _04297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A2 _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ net743 _04991_ net459 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__and3_1
X_06832_ _02935_ _02936_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05705__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__C net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ net217 net2169 net304 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__mux2_1
X_06763_ core.register_file.registers_state\[977\] core.register_file.registers_state\[1009\]
+ net886 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__mux2_1
X_08502_ _04582_ _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05714_ net1057 core.register_file.registers_state\[213\] vssd1 vssd1 vccd1 vccd1
+ _01819_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09482_ _04995_ net323 net263 net1726 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__a22o_1
X_06694_ core.register_file.registers_state\[19\] core.register_file.registers_state\[51\]
+ core.register_file.registers_state\[147\] core.register_file.registers_state\[179\]
+ net871 net819 vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__mux4_1
XANTENNA__06239__C net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08433_ core.pc.current_pc\[18\] _04502_ core.pc.current_pc\[19\] vssd1 vssd1 vccd1
+ vccd1 _04521_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05645_ net949 core.register_file.registers_state\[886\] net764 vssd1 vssd1 vccd1
+ vccd1 _01750_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05703__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08364_ net209 _04458_ net597 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__o21ai_1
X_05576_ net922 _01677_ _01678_ _01680_ net932 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_138_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09445__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07315_ _03418_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__nand2_1
XANTENNA__09996__B2 _05098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08295_ core.pc.current_pc\[7\] _03172_ net577 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1157_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07246_ net773 _03330_ _03337_ _03350_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_95_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07177_ core.register_file.registers_state\[867\] core.register_file.registers_state\[835\]
+ net855 vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__mux2_1
XANTENNA__09566__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout203_X net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06128_ core.register_file.registers_state\[8\] core.register_file.registers_state\[40\]
+ net700 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XANTENNA__08420__A1 _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout784_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06059_ net651 _02161_ _02163_ net958 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1112_X net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1308 net1312 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__clkbuf_2
Xfanout310 _05063_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_4
Xfanout332 _05047_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_4
Xfanout343 _05027_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout951_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 net356 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_4
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_8
Xfanout376 net377 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08723__A2 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09818_ _04884_ net2222 net381 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
Xfanout387 net389 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_4
Xfanout398 net404 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06734__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__B1 _03937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_clk_X clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _04967_ net295 net258 net1750 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__a22o_1
XANTENNA__05942__C1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09684__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08926__A _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11711_ clknet_leaf_52_clk net1526 net1303 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08239__A1 _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11642_ clknet_leaf_52_clk _01154_ net1303 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09436__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05350__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10046__B2 core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09987__B2 _02451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11573_ clknet_leaf_27_clk _01085_ net1197 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07998__B1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_1
XFILLER_0_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10524_ clknet_leaf_32_clk _00036_ net1207 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[28\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05473__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05473__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06670__B1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ net1355 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10386_ net1418 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06973__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08175__B1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09911__A1 core.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ clknet_leaf_14_clk _00519_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[479\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05528__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06725__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06725__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_101_clk_X clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09675__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05430_ net1047 core.register_file.registers_state\[190\] net674 core.register_file.registers_state\[158\]
+ net639 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09003__Y _04975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05260__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05361_ net785 _01464_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07100_ _03200_ _03203_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__or2_1
X_08080_ _04025_ _04071_ _04180_ _04184_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05292_ core.decoder.inst\[14\] _01397_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_133_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07031_ net1103 core.register_file.registers_state\[840\] core.register_file.registers_state\[872\]
+ net838 net981 vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__o221a_1
XANTENNA__06661__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07187__A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05419__B net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ net611 _04662_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07933_ _03927_ _04037_ net531 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08510__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07864_ _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06716__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09603_ net2236 net394 _05067_ net1000 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__a22o_1
X_06815_ net1091 core.register_file.registers_state\[333\] core.register_file.registers_state\[365\]
+ net831 net978 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__o221a_1
X_07795_ _02598_ _03536_ net580 vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06811__S1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout365_A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09534_ net207 net2395 net304 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06746_ net1111 core.register_file.registers_state\[337\] core.register_file.registers_state\[369\]
+ net857 net983 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09666__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09465_ _04704_ net2036 net263 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout532_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06677_ net551 _02781_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06575__S0 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08416_ _01958_ _04504_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__nand2_1
X_05628_ core.register_file.registers_state\[23\] net671 net653 _01732_ vssd1 vssd1
+ vccd1 vccd1 _01733_ sky130_fd_sc_hd__a211o_1
XANTENNA__06266__A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ net1842 net329 net321 _04876_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07429__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ _02117_ _04442_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05559_ net584 _01646_ _01663_ _01634_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout1062_X net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08278_ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__inv_2
XANTENNA__08481__A _01710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06247__A3 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout999_A _01368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07229_ net989 core.register_file.registers_state\[705\] net875 core.register_file.registers_state\[737\]
+ net809 vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07097__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ net1126 net1444 net911 _05228_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_37_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09197__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10235__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10200__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net129 net916 net906 net1581 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a22o_1
XANTENNA__05329__B core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 net1106 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_4
Xfanout1116 net1117 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_4
Xfanout1127 _01379_ vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1138 net1139 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08157__B1 _02017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10251__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06707__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11135__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09657__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_70_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07132__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05694__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ clknet_leaf_72_clk _01137_ net1269 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08093__C1 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ clknet_leaf_26_clk _01068_ net1191 vssd1 vssd1 vccd1 vccd1 core.control_logic.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire552 _02686_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_4
XFILLER_0_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05446__A1 core.decoder.inst\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10507_ clknet_leaf_45_clk _00019_ net1288 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06643__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11487_ clknet_leaf_62_clk _00999_ net1242 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[959\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09188__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10438_ net1377 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07199__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ _05121_ net1608 net232 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__mux2_1
XANTENNA__06946__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09426__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08148__B1 _03950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_23_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07454__B net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05255__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05906__C1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ net1106 core.register_file.registers_state\[182\] net851 core.register_file.registers_state\[150\]
+ net810 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07580_ _02384_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__nor2_4
XANTENNA__05382__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09648__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10258__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06531_ core.register_file.registers_state\[28\] core.register_file.registers_state\[60\]
+ core.register_file.registers_state\[156\] core.register_file.registers_state\[188\]
+ net873 net822 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux4_1
XANTENNA__10502__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09250_ core.register_file.registers_state\[316\] net475 net545 net560 vssd1 vssd1
+ vccd1 vccd1 _05041_ sky130_fd_sc_hd__o211a_1
X_06462_ net1037 net747 core.register_file.registers_state\[536\] vssd1 vssd1 vccd1
+ vccd1 _02567_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06331__C1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ net527 _03965_ _04299_ _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__o31a_2
XFILLER_0_111_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05685__A1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05413_ net1047 core.register_file.registers_state\[734\] core.register_file.registers_state\[766\]
+ net674 net654 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__o221a_1
X_06393_ _02493_ _02497_ net657 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
X_09181_ _04967_ net359 net425 net2111 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05780__S1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05344_ wb.curr_state\[0\] _01451_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__nand2_1
X_08132_ net478 _03760_ _03763_ net491 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08623__A1 core.IO_mod.input_reg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09820__A0 _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload52_A clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ _03868_ _03869_ _04086_ _03892_ net482 net492 vssd1 vssd1 vccd1 vccd1 _04168_
+ sky130_fd_sc_hd__mux4_2
X_05275_ core.control_logic.instruction\[1\] core.control_logic.instruction\[0\] core.control_logic.instruction\[2\]
+ core.control_logic.instruction\[3\] vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_77_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09179__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07014_ net785 _03117_ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10055__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10194__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1022_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08965_ _04855_ net601 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout482_A _02516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ net1003 _02016_ _02962_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_23_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08896_ _04730_ net737 vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__and2_1
XANTENNA__09887__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__X _04037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09351__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ _01612_ _02660_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ _03697_ _03867_ _03878_ _03882_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o211a_2
XANTENNA__09639__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05912__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07380__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ _04802_ net397 net307 net1949 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09103__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06729_ net1110 core.register_file.registers_state\[594\] core.register_file.registers_state\[626\]
+ net860 net813 vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout914_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1277_X net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09448_ _04930_ net318 net312 net2049 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__a22o_1
XANTENNA__06322__C1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05676__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06873__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ net1710 net327 net315 _04786_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__a22o_1
XANTENNA__08923__B net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05771__S1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ clknet_leaf_64_clk _00922_ net1249 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[882\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09811__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05428__A1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ clknet_leaf_2_clk _00853_ net1139 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[813\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11272_ clknet_leaf_14_clk _00784_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[744\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10223_ net72 net920 vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__and2_1
XANTENNA__06389__C1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10185__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07555__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _03811_ _05190_ net255 vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__or3b_1
XFILLER_0_24_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09590__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05600__B2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10085_ net1602 net517 net472 _05150_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__a22o_1
Xhold7 core.register_file.registers_state\[929\] vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08145__A3 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10987_ clknet_leaf_111_clk _00499_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[459\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05522__B _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05667__A1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11608_ clknet_leaf_27_clk _01120_ net1197 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09802__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09010__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11539_ clknet_leaf_11_clk _01051_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1011\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08081__A2 _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold407 core.register_file.registers_state\[529\] vssd1 vssd1 vccd1 vccd1 net1726
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold418 core.register_file.registers_state\[671\] vssd1 vssd1 vccd1 vccd1 net1737
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11236__RESET_B net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold429 core.register_file.registers_state\[902\] vssd1 vssd1 vccd1 vccd1 net1748
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10176__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout909 _05205_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09581__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 core.register_file.registers_state\[585\] vssd1 vssd1 vccd1 vccd1 net2426
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05256__Y _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08750_ net2205 net469 net438 _04807_ vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_124_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 core.register_file.registers_state\[138\] vssd1 vssd1 vccd1 vccd1 net2437
+ sky130_fd_sc_hd__dlygate4sd3_1
X_05962_ core.register_file.registers_state\[557\] net666 vssd1 vssd1 vccd1 vccd1
+ _02067_ sky130_fd_sc_hd__or2_1
Xhold1129 core.register_file.registers_state\[320\] vssd1 vssd1 vccd1 vccd1 net2448
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ net451 _03446_ net443 net505 vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__a31o_1
XANTENNA__09333__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08681_ core.IO_mod.input_reg\[7\] net252 net725 vssd1 vssd1 vccd1 vccd1 _04749_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05893_ core.register_file.registers_state\[175\] net681 net658 _01997_ vssd1 vssd1
+ vccd1 vccd1 _01998_ sky130_fd_sc_hd__o211a_1
X_07632_ _03611_ _03610_ net255 vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08296__A core.decoder.inst\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05713__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07563_ _03660_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09302_ _04917_ net417 net332 net1996 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09679__X _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06514_ net1082 _02618_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_17_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07494_ net791 _03595_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05658__A1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ net559 _04817_ _05032_ net340 net2442 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_118_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06445_ net1063 core.register_file.registers_state\[89\] core.register_file.registers_state\[121\]
+ net690 net649 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_79_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09398__Y _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08743__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09164_ _04936_ net355 net344 net2204 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__a22o_1
X_06376_ core.register_file.registers_state\[866\] core.register_file.registers_state\[834\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XANTENNA__10337__Y _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ net477 _03351_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__nand2_1
X_05327_ _01439_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09095_ net2490 net366 net359 _04806_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1237_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08046_ _02276_ _03172_ net578 vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__o21a_1
X_05258_ net1025 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
Xhold930 core.register_file.registers_state\[324\] vssd1 vssd1 vccd1 vccd1 net2249
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold941 core.register_file.registers_state\[111\] vssd1 vssd1 vccd1 vccd1 net2260
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05830__A1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout697_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold952 core.register_file.registers_state\[36\] vssd1 vssd1 vccd1 vccd1 net2271
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 core.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold974 core.register_file.registers_state\[174\] vssd1 vssd1 vccd1 vccd1 net2293
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10167__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold985 core.register_file.registers_state\[459\] vssd1 vssd1 vccd1 vccd1 net2304
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1025_X net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold996 core.register_file.registers_state\[700\] vssd1 vssd1 vccd1 vccd1 net2315
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09572__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07032__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ net594 _02204_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nor2_4
XFILLER_0_122_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ net571 net214 net738 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_4_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08758__X _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05594__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09324__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ net204 net2523 net371 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10910_ clknet_leaf_95_clk _00422_ net1178 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10698__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ clknet_leaf_46_clk _01359_ net1291 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07886__A2 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06543__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10841_ clknet_leaf_68_clk _00353_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07541__C net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05992__S1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05342__B net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10772_ clknet_leaf_53_clk _00284_ net1304 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05910__X _02015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08653__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09260__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06173__B _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06074__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06074__B2 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07271__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ clknet_leaf_41_clk _00836_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[796\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05821__A1 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11255_ clknet_leaf_22_clk _00767_ net1180 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[727\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10206_ net1128 net1550 net913 _05211_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__a31o_1
XANTENNA__07023__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ clknet_leaf_67_clk _00698_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[658\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07574__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10137_ core.pc.current_pc\[29\] _05183_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09315__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ net2055 net518 _05140_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10330__A0 _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07877__A2 _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05888__A1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05533__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09079__B2 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05820__X _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06230_ net629 _02323_ _02328_ net723 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06161_ net1054 core.register_file.registers_state\[679\] core.register_file.registers_state\[647\]
+ net685 net643 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08850__Y _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06065__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold204 core.CPU_DAT_I\[9\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07747__X _03852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11070__RESET_B net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06092_ net1052 core.register_file.registers_state\[329\] vssd1 vssd1 vccd1 vccd1
+ _02197_ sky130_fd_sc_hd__or2_1
XANTENNA__07262__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold215 _01218_ vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 core.CPU_DAT_I\[27\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 core.register_file.registers_state\[299\] vssd1 vssd1 vccd1 vccd1 net1556
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold248 core.CPU_DAT_I\[30\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ net1122 net2068 net891 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__mux2_1
Xhold259 core.register_file.registers_state\[27\] vssd1 vssd1 vccd1 vccd1 net1578
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10149__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 net707 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_4
Xfanout717 net720 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_6
XFILLER_0_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09851_ _04909_ net390 net268 net2100 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
Xfanout739 net740 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
XANTENNA__10164__A3 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08802_ net1868 net469 net438 _04851_ vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__a22o_1
X_09782_ _04726_ net387 net271 net1794 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__a22o_1
X_06994_ core.register_file.registers_state\[777\] core.register_file.registers_state\[809\]
+ core.register_file.registers_state\[905\] core.register_file.registers_state\[937\]
+ net872 net1074 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06773__C1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10840__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08109__A3 _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ core.IO_mod.input_reg\[15\] net253 vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__and2_1
XANTENNA__09306__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05945_ net633 _02046_ _02049_ net723 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout278_A _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ core.IO_mod.input_reg\[4\] net253 net728 vssd1 vssd1 vccd1 vccd1 _04735_
+ sky130_fd_sc_hd__a21oi_1
X_05876_ core.register_file.registers_state\[977\] core.register_file.registers_state\[1009\]
+ net711 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__mux2_1
XANTENNA__07412__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07615_ net497 _03719_ _03718_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08595_ core.decoder.inst\[8\] _04656_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__or2_4
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1187_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07546_ net507 _03646_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nor2_1
XANTENNA__06826__X _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08754__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06828__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07477_ net582 _03566_ _03580_ _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a31oi_4
XANTENNA_fanout612_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11158__RESET_B net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ _04732_ net421 net342 net1746 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__a22o_1
XANTENNA__11346__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06428_ net555 _01745_ _01780_ _01711_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09147_ _04902_ net359 net346 net2219 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06359_ _02460_ _02463_ net630 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_40_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1142_X net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09793__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ net2499 net365 net360 _04707_ vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout981_A _01370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11496__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06151__S1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08029_ _04083_ _04133_ net492 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06280__Y _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold760 core.register_file.registers_state\[450\] vssd1 vssd1 vccd1 vccd1 net2079
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold771 core.IO_mod.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold782 core.register_file.registers_state\[481\] vssd1 vssd1 vccd1 vccd1 net2101
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11040_ clknet_leaf_59_clk _00552_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[512\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold793 core.register_file.registers_state\[73\] vssd1 vssd1 vccd1 vccd1 net2112
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07536__C net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10243__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07552__B _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10312__A0 _02272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06516__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ clknet_leaf_54_clk _01342_ net1299 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10824_ clknet_leaf_12_clk _00336_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[296\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05640__X _01745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10076__C1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06819__B1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ clknet_leaf_71_clk _00267_ net1272 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[227\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06295__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05499__S net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ clknet_leaf_96_clk _00198_ net1174 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[158\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10713__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11839__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09233__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__Y _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07244__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__A1 _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11307_ clknet_leaf_109_clk _00819_ net1134 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[779\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11238_ clknet_leaf_98_clk _00750_ net1160 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[710\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08744__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11169_ clknet_leaf_102_clk _00681_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[641\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08839__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__A _01583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05730_ core.register_file.registers_state\[532\] net714 net649 _01834_ vssd1 vssd1
+ vccd1 vccd1 _01835_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_19_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05661_ core.register_file.registers_state\[214\] core.register_file.registers_state\[246\]
+ net706 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05956__S1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ _03499_ _03504_ net782 vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__mux2_1
XANTENNA__11369__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ _02053_ _04463_ _04451_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05592_ net1041 core.register_file.registers_state\[187\] vssd1 vssd1 vccd1 vccd1
+ _01697_ sky130_fd_sc_hd__and2_1
XANTENNA__05730__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10067__C1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07331_ net969 _03434_ _03435_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09472__A1 _04975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07262_ _03364_ _03366_ net782 vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07483__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06094__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09001_ net612 net568 _04746_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06213_ net941 core.register_file.registers_state\[37\] net761 vssd1 vssd1 vccd1
+ vccd1 _02318_ sky130_fd_sc_hd__or3_1
X_07193_ net994 core.register_file.registers_state\[706\] net884 core.register_file.registers_state\[738\]
+ net815 vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__a221o_1
XANTENNA__09224__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06038__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06144_ net945 core.register_file.registers_state\[199\] net703 core.register_file.registers_state\[231\]
+ net643 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a221o_1
XANTENNA__09775__A2 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07786__A1 _03890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06075_ net1052 core.register_file.registers_state\[969\] core.register_file.registers_state\[1001\]
+ net678 net1015 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__o221a_1
XANTENNA__05797__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ net1115 _05078_ net375 net2344 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__a22o_1
XANTENNA__09527__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout503 _02454_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_2
Xfanout514 _02422_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout525 _04757_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_4
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout395_A net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 _03622_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_4
X_09834_ _04891_ net1906 net380 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1102_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 net559 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_4
XANTENNA__08749__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06746__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 net570 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06210__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ _04999_ net289 net260 net2392 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__a22o_1
X_06977_ _02176_ _03053_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1210_A core.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08716_ net729 _04096_ _04777_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a22o_1
X_05928_ net945 core.register_file.registers_state\[590\] net705 core.register_file.registers_state\[622\]
+ net657 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a221oi_1
X_09696_ _04800_ net2513 net279 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06269__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09160__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08647_ net570 net436 _04720_ net468 net1564 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05859_ net1060 core.register_file.registers_state\[209\] core.register_file.registers_state\[241\]
+ net689 net661 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ net1122 net895 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07529_ net449 net550 net441 net507 vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__o31a_1
XANTENNA__10736__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09463__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10540_ clknet_leaf_102_clk _00052_ net1162 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08671__C1 _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05485__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09215__A1 _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10471_ net1359 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10886__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09766__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06985__C1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09518__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold590 core.register_file.registers_state\[716\] vssd1 vssd1 vccd1 vccd1 net1909
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07529__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ clknet_leaf_82_clk _00535_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[495\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08659__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06201__A1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05555__A3 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05960__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07162__C1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__Y _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11856_ clknet_leaf_28_clk net52 net1195 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11009__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ clknet_leaf_21_clk _00319_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[279\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11787_ clknet_leaf_30_clk _01291_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06268__A1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ clknet_leaf_71_clk _00250_ net1274 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[210\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07465__B1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05476__C1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06363__S1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08009__A2 _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10669_ clknet_leaf_2_clk _00181_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[141\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07217__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09429__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09757__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08333__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XANTENNA__07457__B net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XANTENNA__10644__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05258__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ core.register_file.registers_state\[780\] core.register_file.registers_state\[812\]
+ net870 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07880_ net529 _03966_ _03967_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a31o_4
XANTENNA__08213__A_N _03964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__C1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07473__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06831_ _02931_ _02934_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05264__Y _01379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ net218 net2508 net303 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__mux2_1
X_06762_ core.register_file.registers_state\[913\] core.register_file.registers_state\[945\]
+ net883 vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__mux2_1
XANTENNA__05951__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ core.pc.current_pc\[24\] core.pc.current_pc\[25\] _04562_ vssd1 vssd1 vccd1
+ vccd1 _04583_ sky130_fd_sc_hd__and3_1
X_05713_ net1056 core.register_file.registers_state\[85\] vssd1 vssd1 vccd1 vccd1
+ _01818_ sky130_fd_sc_hd__or2_1
X_09481_ _04993_ net318 net261 net1592 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__a22o_1
X_06693_ net968 _02793_ _02796_ _02797_ _02788_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08432_ core.pc.current_pc\[18\] core.pc.current_pc\[19\] _04502_ vssd1 vssd1 vccd1
+ vccd1 _04520_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07920__B _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05644_ net1056 core.register_file.registers_state\[982\] core.register_file.registers_state\[1014\]
+ net684 net1019 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05721__A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08363_ core.pc.current_pc\[12\] _04440_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05575_ net937 core.register_file.registers_state\[1019\] net758 _01679_ net1012
+ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_138_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07314_ _02720_ _03414_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nor2_1
XANTENNA__06259__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08294_ core.pc.current_pc\[6\] net599 _04392_ _04394_ vssd1 vssd1 vccd1 vccd1 _00014_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08591__X _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07245_ net777 _03342_ _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_95_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout310_A _05063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1052_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09748__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ core.register_file.registers_state\[803\] core.register_file.registers_state\[771\]
+ net855 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__mux2_1
XANTENNA__06552__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06127_ net960 _02228_ _02231_ net627 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10074__A _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06058_ core.register_file.registers_state\[650\] net669 net636 _02162_ vssd1 vssd1
+ vccd1 vccd1 _02163_ sky130_fd_sc_hd__a211o_1
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_8
Xfanout311 _05058_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_6
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1309 net1310 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08708__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout322 net326 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07654__Y _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout333 _05047_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_6
Xfanout344 _05027_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1105_X net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06719__C1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_4
Xfanout366 _05023_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11534__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout377 net378 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_31_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09817_ net223 net2052 net380 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_4
XANTENNA_fanout944_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 net403 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
XANTENNA__07931__B2 _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _04965_ net294 net258 net1860 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__a22o_1
XANTENNA__09133__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ _04654_ net604 _05062_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or3_4
X_11710_ clknet_leaf_52_clk net1496 net1302 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09845__C_N net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08926__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11641_ clknet_leaf_52_clk _01153_ net1302 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11102__RESET_B net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05350__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09987__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ clknet_leaf_29_clk _01084_ net1195 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08942__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07998__A1 _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ clknet_leaf_33_clk _00035_ net1207 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07558__A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ net1354 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09739__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11064__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08411__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10385_ net1431 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05630__C1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08175__B2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07293__A _03139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09372__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ clknet_leaf_95_clk _00518_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07922__A1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05525__B _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08676__X _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07135__C1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06489__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06489__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09013__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ clknet_leaf_36_clk net65 net1223 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09427__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05360_ net1098 core.register_file.registers_state\[222\] core.register_file.registers_state\[254\]
+ net842 net819 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08852__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05291_ _01366_ net896 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07030_ net1103 core.register_file.registers_state\[968\] core.register_file.registers_state\[1000\]
+ net838 net1070 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__o221a_1
XANTENNA__05464__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06661__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08981_ net2323 net369 _04960_ net437 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__a22o_1
X_07932_ _03969_ _03991_ _04013_ _04011_ net479 net495 vssd1 vssd1 vccd1 vccd1 _04037_
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_71_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09363__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07863_ _03645_ _03675_ net498 vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__mux2_1
XANTENNA__09902__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06177__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10581__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09602_ net743 _04965_ net459 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__and3_1
X_06814_ net1091 core.register_file.registers_state\[461\] core.register_file.registers_state\[493\]
+ net831 net1069 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07794_ _02598_ _03536_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__and2_1
XANTENNA__09115__A0 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ _04882_ _05062_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__or2_1
X_06745_ net1111 core.register_file.registers_state\[465\] core.register_file.registers_state\[497\]
+ net857 net1078 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout358_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05722__Y _01827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07650__B _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _04961_ net319 vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__nand2_2
X_06676_ _01865_ _02780_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08415_ _01958_ _04504_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__or2_1
XANTENNA__05688__C1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06575__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05627_ net1041 core.register_file.registers_state\[55\] net749 vssd1 vssd1 vccd1
+ vccd1 _01732_ sky130_fd_sc_hd__and3_1
XANTENNA__09418__A1 _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ net1769 net327 net317 _04871_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08346_ core.pc.current_pc\[11\] _03052_ net576 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__mux2_1
XANTENNA__10028__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05558_ net717 _01655_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__or3_2
XFILLER_0_62_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08277_ core.decoder.inst\[25\] _01412_ _04377_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a21oi_2
X_05489_ core.register_file.registers_state\[92\] core.register_file.registers_state\[124\]
+ net699 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07228_ net824 _03331_ _03332_ net974 vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__o211a_1
XANTENNA__06652__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06652__B2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06282__A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07159_ _03261_ _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08610__D_N _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ net128 net917 net907 net1479 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_2
XANTENNA__05612__C1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1117 core.decoder.inst\[10\] vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_4
Xfanout1128 _01379_ vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1139 net1140 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08157__B2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09354__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10251__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07365__C1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05915__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07841__A _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07117__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05361__A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11624_ clknet_leaf_71_clk _01136_ net1270 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08672__A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11555_ clknet_leaf_26_clk _01067_ net1208 vssd1 vssd1 vccd1 vccd1 core.control_logic.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire553 _02659_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_4
X_10506_ clknet_leaf_37_clk _00018_ net1222 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05446__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11486_ clknet_leaf_93_clk _00998_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[958\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10437_ net1335 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09707__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09593__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10368_ _05120_ net2059 net232 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__mux2_1
XANTENNA__06920__A _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10299_ net22 net902 net796 net2422 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08148__B2 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10161__B net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07356__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05906__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09648__A1 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05382__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06530_ _02630_ _02632_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06461_ net943 core.register_file.registers_state\[568\] net760 vssd1 vssd1 vccd1
+ vccd1 _02566_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08200_ _03685_ _04169_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05412_ net1048 core.register_file.registers_state\[606\] core.register_file.registers_state\[638\]
+ net679 net640 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__o221a_1
X_09180_ _04965_ net361 net425 net1786 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06882__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06392_ net944 core.register_file.registers_state\[673\] core.register_file.registers_state\[641\]
+ net702 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08582__A core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _04160_ _04210_ net478 vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05343_ core.READ_I core.WRITE_I vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08623__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06095__C1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06634__A1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ _02316_ _03201_ net547 _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05274_ core.control_logic.instruction\[1\] core.control_logic.instruction\[0\] core.control_logic.instruction\[2\]
+ core.control_logic.instruction\[3\] vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_77_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10947__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07013_ net1100 core.register_file.registers_state\[200\] core.register_file.registers_state\[232\]
+ net843 net821 vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__o221a_1
XANTENNA__05842__C1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09584__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06830__A _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06398__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08964_ net2356 net370 _04949_ net439 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1015_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _02016_ _02962_ net578 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06041__S net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ net2412 net369 _04903_ net438 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout475_A _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _03949_ _03950_ net511 vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07777_ net511 _03879_ _03881_ _03658_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__a211o_1
XANTENNA__05373__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05373__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ _04797_ net400 net309 net1851 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a22o_1
X_06728_ net1110 core.register_file.registers_state\[722\] core.register_file.registers_state\[754\]
+ net860 net828 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06277__A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09447_ _04928_ net321 net313 net2156 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06659_ net781 _02755_ _02758_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_42_clk_X clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1172_X net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout907_A _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06873__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ net1870 net328 net320 _04781_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__a22o_1
XANTENNA__11722__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08329_ core.pc.current_pc\[9\] net597 _04418_ _04426_ vssd1 vssd1 vccd1 vccd1 _00017_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09811__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11340_ clknet_leaf_103_clk _00852_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[812\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06443__C net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11271_ clknet_leaf_91_clk _00783_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[743\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10222_ net1127 net1443 net912 _05219_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09575__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06740__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06389__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ _03811_ _05190_ net255 vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07555__B _03659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08003__Y _04108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_A gpio_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ core.pc.current_pc\[13\] _04075_ net590 vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__mux2_1
XANTENNA__07338__C1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 core.register_file.registers_state\[985\] vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08667__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09262__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10986_ clknet_leaf_0_clk _00498_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[458\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06187__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06313__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09498__A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11607_ clknet_leaf_27_clk _01119_ net1204 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09802__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06616__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06616__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09010__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11538_ clknet_leaf_65_clk _01050_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1010\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06353__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold408 core.register_file.registers_state\[270\] vssd1 vssd1 vccd1 vccd1 net1727
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 core.register_file.registers_state\[868\] vssd1 vssd1 vccd1 vccd1 net1738
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11469_ clknet_leaf_1_clk _00981_ net1139 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[941\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08369__A1 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05965__S net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08341__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07041__A1 _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09318__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05961_ _02065_ _02064_ _02060_ _02059_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__o2bb2a_1
Xhold1108 core.register_file.registers_state\[200\] vssd1 vssd1 vccd1 vccd1 net2427
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1119 core.register_file.registers_state\[584\] vssd1 vssd1 vccd1 vccd1 net2438
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07329__C1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ net450 net553 net442 net505 vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__o31a_1
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08680_ net1850 net467 net433 _04748_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_109_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05892_ net1054 core.register_file.registers_state\[143\] vssd1 vssd1 vccd1 vccd1
+ _01997_ sky130_fd_sc_hd__or2_1
XANTENNA__08577__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06001__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07631_ net537 net529 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08296__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07562_ net483 _03661_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_66_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09097__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09301_ _04915_ net417 net331 net2014 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06513_ core.register_file.registers_state\[797\] core.register_file.registers_state\[829\]
+ core.register_file.registers_state\[925\] core.register_file.registers_state\[957\]
+ net868 net1070 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_17_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07493_ net786 _03596_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__or3_1
XFILLER_0_76_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ core.register_file.registers_state\[307\] net475 net545 vssd1 vssd1 vccd1
+ vccd1 _05032_ sky130_fd_sc_hd__o21a_1
X_06444_ core.register_file.registers_state\[25\] net690 net662 _02548_ vssd1 vssd1
+ vccd1 vccd1 _02549_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07420__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08743__C net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ _04934_ net360 net345 net2108 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__a22o_1
X_06375_ core.register_file.registers_state\[802\] core.register_file.registers_state\[770\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout223_A _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08114_ net547 _04218_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__nor2_1
X_05326_ net1315 _01421_ _01438_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__a21o_1
X_09094_ net2203 net363 net353 _04801_ vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05815__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ _02276_ _03172_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06083__A2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05257_ net1068 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_4
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold920 core.register_file.registers_state\[615\] vssd1 vssd1 vccd1 vccd1 net2239
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1132_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold931 core.register_file.registers_state\[231\] vssd1 vssd1 vccd1 vccd1 net2250
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09557__A0 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05875__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold942 core.register_file.registers_state\[737\] vssd1 vssd1 vccd1 vccd1 net2261
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 core.register_file.registers_state\[839\] vssd1 vssd1 vccd1 vccd1 net2272
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 core.register_file.registers_state\[78\] vssd1 vssd1 vccd1 vccd1 net2283
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A _05093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 core.register_file.registers_state\[497\] vssd1 vssd1 vccd1 vccd1 net2294
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold986 core.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold997 core.register_file.registers_state\[118\] vssd1 vssd1 vccd1 vccd1 net2316
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__A _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ net1476 net540 net519 _05098_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09309__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ net214 net738 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11275__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08878_ net741 _04860_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__nor2_1
XANTENNA__07966__S0 _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07829_ _03821_ _03933_ net481 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ clknet_leaf_10_clk _00352_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[312\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09088__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_99_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ clknet_leaf_12_clk _00283_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[243\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06310__A3 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08653__C net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10257__A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06059__C1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09796__B1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08950__A _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11323_ clknet_leaf_23_clk _00835_ net1182 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[795\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05806__C1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07271__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05282__B1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__A0 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_37_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11254_ clknet_leaf_59_clk _00766_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[726\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08014__X _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10205_ net94 net920 vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07023__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05357__Y _01462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11185_ clknet_leaf_81_clk _00697_ net1255 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[657\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10136_ net470 _05185_ _05186_ net515 net1463 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10067_ _04172_ net557 net591 core.pc.current_pc\[6\] net472 vssd1 vssd1 vccd1 vccd1
+ _05140_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11768__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09720__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09079__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10792__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ clknet_leaf_68_clk _00481_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[441\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10094__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06298__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06645__A _02747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09021__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11148__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06160_ core.register_file.registers_state\[551\] core.register_file.registers_state\[519\]
+ net685 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XANTENNA__09787__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08860__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold205 _01210_ vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06091_ core.register_file.registers_state\[265\] core.register_file.registers_state\[297\]
+ core.register_file.registers_state\[393\] core.register_file.registers_state\[425\]
+ net699 net1015 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux4_1
Xhold216 net147 vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _01228_ vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold238 core.register_file.registers_state\[558\] vssd1 vssd1 vccd1 vccd1 net1557
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _01231_ vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07476__A core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06470__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09850_ _04907_ net387 net267 net1738 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__a22o_1
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_4
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_8
Xfanout729 net730 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08762__B2 _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ net571 net609 net211 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__and3_2
X_06993_ _03094_ _03097_ net772 _03092_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a211o_1
XANTENNA__05576__A1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ net569 _04720_ net390 net272 net1522 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08732_ net729 _04028_ _04757_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__a21oi_1
X_05944_ _02047_ _02048_ net963 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08514__A1 _03475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07415__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ core.IO_mod.data_from_mem\[4\] net248 vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nand2_2
X_05875_ core.register_file.registers_state\[849\] core.register_file.registers_state\[881\]
+ net709 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ net449 _03382_ net441 vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__or3_1
X_08594_ core.decoder.inst\[8\] _04656_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__nor2_2
XFILLER_0_7_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07545_ _03639_ _03649_ net496 vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__mux2_2
XFILLER_0_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout340_A _05031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08754__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06289__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ core.decoder.inst\[31\] net584 vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06555__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09490__A2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06427_ _01866_ _02531_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__nor2_1
X_09215_ _04726_ net421 net341 net1806 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__a22o_1
XANTENNA__05500__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05500__B2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout226_X net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07938__X _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09146_ _04900_ net357 net345 net2007 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__a22o_1
X_06358_ net623 _02461_ _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_40_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10515__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__C1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05309_ net1129 net1691 _01421_ _01423_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07253__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ net567 _04714_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__nor2_1
XANTENNA__07253__B2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06289_ net953 core.register_file.registers_state\[67\] net711 core.register_file.registers_state\[99\]
+ net661 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08028_ _04099_ _04132_ net478 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold750 core.register_file.registers_state\[624\] vssd1 vssd1 vccd1 vccd1 net2069
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout974_A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold761 core.register_file.registers_state\[238\] vssd1 vssd1 vccd1 vccd1 net2080
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold772 core.register_file.registers_state\[636\] vssd1 vssd1 vccd1 vccd1 net2091
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07005__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold783 core.register_file.registers_state\[647\] vssd1 vssd1 vccd1 vccd1 net2102
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 core.register_file.registers_state\[241\] vssd1 vssd1 vccd1 vccd1 net2113
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10665__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05567__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ net1129 core.WRITE_I _01423_ _01427_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__B net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__B _03937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__A2 _03412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11872_ clknet_leaf_50_clk _01341_ net1310 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08945__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09540__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08269__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10823_ clknet_leaf_92_clk _00335_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[295\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10076__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06819__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754_ clknet_leaf_77_clk _00266_ net1258 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[226\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09481__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07492__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685_ clknet_leaf_17_clk _00197_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[157\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07492__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09769__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09233__A2 _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07244__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07795__A2 _03536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11306_ clknet_leaf_1_clk _00818_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[778\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11237_ clknet_leaf_88_clk _00749_ net1229 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[709\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09941__A0 core.decoder.inst\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ clknet_leaf_59_clk _00680_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[640\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06755__B1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08839__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ net1124 core.pc.current_pc\[25\] core.pc.current_pc\[26\] vssd1 vssd1 vccd1
+ vccd1 _05172_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07743__B _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06850__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ clknet_leaf_19_clk _00611_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[571\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09016__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05660_ core.register_file.registers_state\[150\] core.register_file.registers_state\[182\]
+ net706 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__mux2_1
XANTENNA__05715__D1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05591_ core.register_file.registers_state\[27\] net671 net653 _01695_ vssd1 vssd1
+ vccd1 vccd1 _01696_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_109_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10067__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07330_ net1095 core.register_file.registers_state\[603\] core.register_file.registers_state\[635\]
+ net837 net803 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09472__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10538__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07261_ net1090 _03362_ _03365_ net983 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06286__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07483__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08680__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ net612 _04746_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__and2_1
X_06212_ net1047 core.register_file.registers_state\[133\] net674 core.register_file.registers_state\[165\]
+ net655 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__o221a_1
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06691__C1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07192_ net995 core.register_file.registers_state\[578\] net883 core.register_file.registers_state\[610\]
+ net827 vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06143_ net948 core.register_file.registers_state\[71\] net706 core.register_file.registers_state\[103\]
+ net659 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07477__Y _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__A3 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06074_ net1051 core.register_file.registers_state\[841\] core.register_file.registers_state\[873\]
+ net678 net925 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_93_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09902_ _05007_ net384 net375 net1836 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout504 _02453_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
Xfanout515 _05126_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07538__A2 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__A0 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout526 _04756_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_4
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout537 net539 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
X_09833_ net214 net1896 net381 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
Xfanout548 _03621_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_4
XANTENNA__05549__A1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06746__B1 core.register_file.registers_state\[369\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net562 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_4
XANTENNA__08749__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06210__A2 _02314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _04997_ net296 net258 net1699 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06976_ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__inv_2
XANTENNA__07145__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05454__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08715_ core.IO_mod.input_reg\[12\] net253 net730 vssd1 vssd1 vccd1 vccd1 _04778_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05927_ net945 core.register_file.registers_state\[718\] vssd1 vssd1 vccd1 vccd1
+ _02032_ sky130_fd_sc_hd__nand2_1
X_09695_ net219 net2269 net280 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout555_A _01506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1297_A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08646_ net610 net226 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__and2_2
X_05858_ net1060 core.register_file.registers_state\[81\] core.register_file.registers_state\[113\]
+ net689 net647 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__o221a_1
XANTENNA__07171__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05789_ net582 _01868_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout722_A _01511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ net1116 net895 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1085_X net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07528_ net450 _02840_ net442 net502 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o31a_1
XANTENNA__06285__A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11463__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07474__A1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05620__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07459_ core.register_file.registers_state\[863\] net707 _03552_ vssd1 vssd1 vccd1
+ vccd1 _03564_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10470_ net1325 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09215__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09129_ _04810_ net2502 net349 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07777__A2 _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05788__B2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 core.register_file.registers_state\[901\] vssd1 vssd1 vccd1 vccd1 net1899
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07529__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 core.register_file.registers_state\[633\] vssd1 vssd1 vccd1 vccd1 net1910
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09923__A0 core.decoder.inst\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09535__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ clknet_leaf_88_clk _00534_ net1229 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[494\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08659__B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10270__A core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05364__A core.decoder.inst\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07701__A2 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09270__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11855_ clknet_leaf_22_clk net51 net1181 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10806_ clknet_leaf_60_clk _00318_ net1284 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[278\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06195__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11786_ clknet_leaf_24_clk _01290_ net1185 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09454__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06899__S0 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737_ clknet_leaf_72_clk _00249_ net1269 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[209\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11049__RESET_B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10668_ clknet_leaf_102_clk _00180_ net1162 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[140\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09206__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07217__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10599_ clknet_leaf_63_clk _00111_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[71\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_131_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08178__C1 _04282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07076__S0 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06830_ _02931_ _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nor2_1
XANTENNA__11336__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06761_ _02862_ _02863_ _02865_ _02864_ net792 net812 vssd1 vssd1 vccd1 vccd1 _02866_
+ sky130_fd_sc_hd__mux4_1
X_08500_ net1124 _04562_ core.pc.current_pc\[25\] vssd1 vssd1 vccd1 vccd1 _04582_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05712_ net949 core.register_file.registers_state\[117\] net763 vssd1 vssd1 vccd1
+ vccd1 _01817_ sky130_fd_sc_hd__or3_1
X_09480_ _04991_ net323 net263 net1803 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a22o_1
X_06692_ net970 _02789_ _02790_ net1066 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_86_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08431_ core.pc.current_pc\[18\] net597 _04517_ _04519_ vssd1 vssd1 vccd1 vccd1 _00026_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05643_ core.register_file.registers_state\[790\] core.register_file.registers_state\[822\]
+ core.register_file.registers_state\[918\] core.register_file.registers_state\[950\]
+ net706 net1019 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__mux4_1
XANTENNA_wire409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11819__RESET_B net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11486__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05703__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05703__B2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05280__Y _01395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08362_ net230 _04455_ _04456_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05574_ net1042 core.register_file.registers_state\[987\] vssd1 vssd1 vccd1 vccd1
+ _01679_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09445__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07313_ _02690_ _02691_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_138_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08293_ net209 _04393_ net599 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_99_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05467__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06664__C1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ net777 _03345_ _03348_ net773 vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11401__RESET_B net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07175_ net995 core.register_file.registers_state\[707\] net887 core.register_file.registers_state\[739\]
+ net983 vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout303_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1045_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06126_ _02229_ _02230_ net1027 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06044__S net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10074__B net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06057_ net1037 core.register_file.registers_state\[682\] vssd1 vssd1 vccd1 vccd1
+ _02162_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1212_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 net302 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout312 _05058_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09905__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout323 net325 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout334 _05047_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout672_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _05027_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_6
Xfanout356 net362 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
Xfanout367 _04898_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_8
X_09816_ net224 net2123 net380 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
XANTENNA__10090__A _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout378 _05089_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout389 net390 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_2
XANTENNA__07931__A2 _03920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _04963_ net292 net259 net1733 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__a22o_1
X_06959_ core.register_file.registers_state\[1002\] core.register_file.registers_state\[970\]
+ net832 vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XANTENNA__05942__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10154__C_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09678_ net607 net241 net291 net283 net1784 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07695__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ _04702_ net244 vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__nand2_8
XFILLER_0_90_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11640_ clknet_leaf_54_clk _01152_ net1299 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09436__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11571_ clknet_leaf_25_clk _01083_ net1191 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08942__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10522_ clknet_leaf_35_clk _00034_ net1220 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11209__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10453_ net1404 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10384_ net1438 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input66_A gpio_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07845__Y _03950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09265__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11005_ clknet_leaf_18_clk _00517_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[477\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06186__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 _01457_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_2
XFILLER_0_137_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07580__Y _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07135__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08883__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11838_ clknet_leaf_22_clk net64 net1181 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05676__B1_N _01779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11769_ clknet_leaf_24_clk _01273_ net1196 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08852__B _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07749__A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05290_ net1123 _01399_ _01403_ _01404_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__or4b_1
XANTENNA__06110__A1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10865__RESET_B net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ net567 net241 net736 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__and3_2
X_07931_ _03774_ _03920_ _03937_ _03798_ _04035_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_71_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10726__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09363__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ _03414_ _03418_ _03965_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_127_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09601_ net999 _04964_ net461 net393 net2164 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06813_ core.register_file.registers_state\[269\] core.register_file.registers_state\[301\]
+ core.register_file.registers_state\[397\] core.register_file.registers_state\[429\]
+ net865 net1069 vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux4_1
X_07793_ net488 _03897_ _03896_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a21o_1
XANTENNA__05924__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09532_ _04881_ net399 net308 net1877 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06744_ core.register_file.registers_state\[273\] core.register_file.registers_state\[305\]
+ core.register_file.registers_state\[401\] core.register_file.registers_state\[433\]
+ net885 net1078 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_84_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09666__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05732__A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ net537 _02531_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__nand2_1
XANTENNA__07221__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08874__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ net241 net735 net319 net312 net1845 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08414_ core.pc.current_pc\[17\] _02873_ net576 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__mux2_1
XANTENNA__06885__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05626_ net1041 core.register_file.registers_state\[183\] net671 core.register_file.registers_state\[151\]
+ net638 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09394_ net1816 net328 net322 _04866_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07429__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08345_ core.pc.current_pc\[11\] _04427_ net229 vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__o21ai_1
X_05557_ net1026 _01656_ _01661_ net1004 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout420_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1162_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06637__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09210__Y _05029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08276_ core.decoder.inst\[25\] net734 _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06101__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05488_ core.register_file.registers_state\[28\] core.register_file.registers_state\[60\]
+ net700 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07227_ net1107 core.register_file.registers_state\[673\] core.register_file.registers_state\[641\]
+ net849 net809 vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06282__B _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07158_ _02384_ _03262_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06109_ net1037 net749 core.register_file.registers_state\[776\] vssd1 vssd1 vccd1
+ vccd1 _02214_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout887_A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07062__C1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10200__A3 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07089_ core.register_file.registers_state\[294\] core.register_file.registers_state\[262\]
+ core.register_file.registers_state\[422\] core.register_file.registers_state\[390\]
+ net842 net1073 vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__mux4_1
XANTENNA__05612__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1107 core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_4
Xfanout1129 _01367_ vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__buf_2
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08157__A2 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09354__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__C_N net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09813__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05376__C1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07460__S0 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07841__B _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07117__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09657__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11394__RESET_B net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__A0 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06876__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08953__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11031__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11623_ clknet_leaf_71_clk _01135_ net1270 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08672__B _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_13_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07569__A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08093__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06628__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11554_ clknet_leaf_26_clk _01066_ net1203 vssd1 vssd1 vccd1 vccd1 core.control_logic.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08017__X _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10505_ clknet_leaf_37_clk _00017_ net1222 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11485_ clknet_leaf_19_clk _00997_ net1190 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[957\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10436_ net1434 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10367_ _05119_ net1890 net235 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__mux2_1
X_10298_ net21 net902 net796 net2134 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_89_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05906__A1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05367__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07108__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09648__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05552__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire221_A _04790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07659__A1 _03763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09024__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10258__A3 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06460_ net1035 net747 core.register_file.registers_state\[920\] vssd1 vssd1 vccd1
+ vccd1 _02565_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06331__A1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05411_ net1008 net747 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__nand2_4
XFILLER_0_29_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06391_ _02494_ _02495_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05685__A3 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08582__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08130_ _03798_ _03890_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05342_ net1 net910 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07479__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08061_ _01365_ _02315_ _03200_ _04165_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a31o_1
XANTENNA__07831__A1 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05273_ net1123 core.control_logic.instruction\[5\] core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_71_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07012_ net1100 core.register_file.registers_state\[72\] core.register_file.registers_state\[104\]
+ net843 net806 vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_77_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09584__A1 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07418__S net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ net571 net211 net738 vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__and3_2
XANTENNA__09336__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ _02016_ _02962_ net548 _01988_ net901 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__a32o_1
X_08894_ net572 net225 net737 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__and3_2
XANTENNA__09887__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__A1 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ _03763_ _03825_ _03887_ net491 vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o22ai_4
XANTENNA__11834__RESET_B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A _04898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ net514 _03880_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__nor2_1
XANTENNA__09639__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07006__X _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ net570 _04791_ net400 net309 net1557 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a32o_1
XANTENNA__11054__CLK clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06727_ net1088 _02828_ _02831_ net1067 vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06277__B _02347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A _01521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ _04926_ net321 net313 net2002 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _02759_ _02760_ _02761_ _02762_ net793 net813 vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06322__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08773__A _04670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05609_ net1043 net749 core.register_file.registers_state\[535\] vssd1 vssd1 vccd1
+ vccd1 _01714_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ net1822 net327 net315 _04776_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout802_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06589_ _02692_ _02693_ net794 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_62_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08328_ net229 _04424_ _04425_ net597 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__o31ai_1
XANTENNA__08075__A1 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07822__A1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ _04361_ _04362_ net598 vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11270_ clknet_leaf_98_clk _00782_ net1160 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[742\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10221_ net71 net920 vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__and2_1
XANTENNA__06389__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10185__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ net588 _05198_ _05199_ net470 vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__o31a_1
XFILLER_0_101_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06232__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10083_ net472 _05148_ _05149_ net517 net1443 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__a32o_1
XANTENNA__08948__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09543__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 core.register_file.registers_state\[939\] vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06010__B1 core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08667__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05372__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08838__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ clknet_leaf_38_clk _00497_ net1217 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09779__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11547__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06313__A1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05667__A3 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__B net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08066__A1 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11606_ clknet_leaf_25_clk _01118_ net1193 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06077__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07274__C1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11537_ clknet_leaf_90_clk _01049_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1009\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09010__C _04888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold409 core.register_file.registers_state\[273\] vssd1 vssd1 vccd1 vccd1 net1728
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11468_ clknet_leaf_103_clk _00980_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[940\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_111_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07026__C1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ net1375 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10176__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ clknet_leaf_65_clk _00911_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[871\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07238__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09019__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05960_ net958 _02061_ net628 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 core.register_file.registers_state\[221\] vssd1 vssd1 vccd1 vccd1 net2428
+ sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_124_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11077__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05891_ core.register_file.registers_state\[47\] core.register_file.registers_state\[15\]
+ net681 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08577__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ _03608_ _03609_ net255 vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__mux2_1
XANTENNA__11245__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07561_ net476 _03662_ _03663_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_66_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09300_ _04913_ net420 net333 net1809 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__a22o_1
X_06512_ _02613_ _02616_ net771 _02611_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_17_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07492_ net1104 core.register_file.registers_state\[223\] core.register_file.registers_state\[255\]
+ net850 net825 vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__o221a_1
XANTENNA__10100__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ _04812_ net421 net342 net1732 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__a22o_1
X_06443_ net1063 core.register_file.registers_state\[57\] net755 vssd1 vssd1 vccd1
+ vccd1 _02548_ sky130_fd_sc_hd__and3_1
XANTENNA__10914__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06374_ core.register_file.registers_state\[930\] core.register_file.registers_state\[898\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
X_09162_ _04932_ net359 net346 net2113 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10880__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05325_ _01422_ _01428_ _01438_ net1473 _01367_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a32o_1
X_08113_ net482 _03352_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07265__C1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ net2262 net365 net357 _04796_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload104_A clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout216_A _04810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net532 _04148_ _03686_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__a21o_1
X_05256_ net1084 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkinv_4
Xhold910 core.register_file.registers_state\[106\] vssd1 vssd1 vccd1 vccd1 net2229
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 core.register_file.registers_state\[335\] vssd1 vssd1 vccd1 vccd1 net2240
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold932 core.register_file.registers_state\[482\] vssd1 vssd1 vccd1 vccd1 net2251
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07017__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold943 core.register_file.registers_state\[175\] vssd1 vssd1 vccd1 vccd1 net2262
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07656__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold954 core.register_file.registers_state\[871\] vssd1 vssd1 vccd1 vccd1 net2273
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1125_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 core.register_file.registers_state\[685\] vssd1 vssd1 vccd1 vccd1 net2284
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10167__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08765__C1 _04819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 core.register_file.registers_state\[419\] vssd1 vssd1 vccd1 vccd1 net2295
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 core.register_file.registers_state\[134\] vssd1 vssd1 vccd1 vccd1 net2306
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 core.register_file.registers_state\[792\] vssd1 vssd1 vccd1 vccd1 net2317
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ net594 net536 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout585_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08946_ net2429 net367 _04937_ net433 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05891__S net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _04893_ net1959 net371 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout752_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07828_ _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__inv_2
XANTENNA__06543__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08605__C_N _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06543__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07759_ net487 _03764_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1282_X net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09599__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ clknet_leaf_69_clk _00282_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[242\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09493__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09429_ net2160 net243 net406 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05503__C1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08048__A1 _03730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__B2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09245__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08008__A _02206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10257__B net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08950__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07847__A _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09538__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ clknet_leaf_8_clk _00834_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[794\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08442__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05282__B2 _01395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07566__B _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11253_ clknet_leaf_63_clk _00765_ net1249 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[725\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11497__SET_B net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10158__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ net1128 net1599 net913 _05210_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11184_ clknet_leaf_104_clk _00696_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[656\]
+ sky130_fd_sc_hd__dfrtp_1
X_10135_ net588 _05181_ _05182_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nand3_1
XANTENNA__06897__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08678__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ net473 _05138_ _05139_ net518 net1655 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__a32o_1
XANTENNA__08030__X _04135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10937__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09484__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10968_ clknet_leaf_10_clk _00480_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[440\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10094__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ clknet_leaf_12_clk _00411_ net1172 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[371\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09021__B _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09236__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08860__B _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06090_ _02191_ _02192_ _02193_ _02194_ net622 net641 vssd1 vssd1 vccd1 vccd1 _02195_
+ sky130_fd_sc_hd__mux4_1
Xhold206 core.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 net201 vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 core.register_file.registers_state\[921\] vssd1 vssd1 vccd1 vccd1 net1547
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07476__B net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 net179 vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08747__C1 _04804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08211__A1 _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 net716 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_2
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout719 net720 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_6
XANTENNA__06222__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08800_ net609 _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__and2_1
XANTENNA__08762__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09780_ net571 _04707_ net388 net271 net1675 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__a32o_1
X_06992_ net971 _03095_ _03096_ net780 vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__o31a_1
XANTENNA__06773__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08588__A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07970__B1 _04073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__B2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09036__X _04997_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ net569 net436 _04791_ net468 net1570 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__a32o_1
X_05943_ net945 core.register_file.registers_state\[462\] net705 core.register_file.registers_state\[494\]
+ net927 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05981__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1290 net1291 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__clkbuf_4
X_08662_ net729 _04255_ _04718_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a21o_1
XANTENNA__06525__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05874_ core.register_file.registers_state\[785\] core.register_file.registers_state\[817\]
+ net711 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
XANTENNA__07722__B1 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08100__B _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09911__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ _03351_ _03631_ net504 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__o21a_1
X_08593_ _04660_ _04663_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and2_2
XANTENNA__08594__Y _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07544_ net479 _03648_ _03644_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09475__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06836__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06289__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07486__C1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07475_ net632 _03579_ _03574_ net722 vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__a211o_2
XFILLER_0_130_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout333_A _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1075_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ net570 _04720_ net419 net341 net1739 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06426_ _02526_ _02530_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09227__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09145_ _04705_ net738 net360 net345 net2041 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout500_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06357_ net952 core.register_file.registers_state\[194\] net710 core.register_file.registers_state\[226\]
+ net646 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1242_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05308_ net1315 core.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08262__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06288_ net953 core.register_file.registers_state\[195\] net714 core.register_file.registers_state\[227\]
+ net649 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09076_ _04714_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08027_ net500 _03703_ _03755_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_57_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__A _04278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 net162 vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 core.register_file.registers_state\[655\] vssd1 vssd1 vccd1 vccd1 net2070
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 core.register_file.registers_state\[329\] vssd1 vssd1 vccd1 vccd1 net2081
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold773 core.IO_mod.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 core.register_file.registers_state\[673\] vssd1 vssd1 vccd1 vccd1 net2103
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold795 core.BUSY_O vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__Y _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout967_A _01372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__A2 _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09978_ net1129 core.READ_I _01428_ _01439_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__a22o_1
X_08929_ net220 net739 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06516__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06516__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09821__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05724__C1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ clknet_leaf_72_clk _01340_ net1271 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10822_ clknet_leaf_100_clk _00334_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[294\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09466__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07341__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10076__A1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05650__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10753_ clknet_leaf_82_clk _00265_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[225\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09218__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06295__A3 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ clknet_leaf_40_clk _00196_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07229__C1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09268__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06452__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ clknet_leaf_16_clk _00817_ net1211 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[777\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11735__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ clknet_leaf_75_clk _00748_ net1257 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[708\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10000__A1 core.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__Y _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__B2 _05100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11167_ clknet_leaf_40_clk _00679_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[639\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06755__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _03946_ _05170_ _05092_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_106_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06850__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11098_ clknet_leaf_9_clk _00610_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[570\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10049_ core.pc.current_pc\[0\] net588 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__or2_1
XANTENNA__09016__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07704__B1 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11115__CLK clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05590_ net1042 core.register_file.registers_state\[59\] net749 vssd1 vssd1 vccd1
+ vccd1 _01695_ sky130_fd_sc_hd__and3_1
XANTENNA__09457__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05730__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10067__A1 _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05560__A core.decoder.inst\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07260_ net996 core.register_file.registers_state\[832\] net888 core.register_file.registers_state\[864\]
+ net977 vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09209__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06211_ net585 _02296_ _02313_ _02278_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07191_ net995 core.register_file.registers_state\[834\] net883 core.register_file.registers_state\[866\]
+ net1078 vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_83_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09224__A3 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05559__X _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06142_ _02244_ _02246_ net618 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__o21a_1
XANTENNA__07487__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05278__Y _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06073_ net1028 _02177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05797__A2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__X _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09901_ net1120 _05077_ net377 net1679 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 _02453_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08196__B1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout516 _05126_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_2
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_4
XANTENNA__09932__A1 core.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ net215 net2365 net382 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06746__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06746__B2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08749__C net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _04995_ net294 net258 net1760 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__a22o_1
X_06975_ net767 _03067_ _03078_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout283_A _05081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_21_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ core.IO_mod.data_from_mem\[12\] net248 vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_33_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09696__A0 _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05926_ core.register_file.registers_state\[750\] net705 vssd1 vssd1 vccd1 vccd1
+ _02031_ sky130_fd_sc_hd__nand2_1
X_09694_ net220 net2310 net280 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09160__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ net728 _04229_ _04716_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_94_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout450_A _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05857_ _01959_ _01961_ net623 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a21o_1
XANTENNA__07171__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ net896 _04650_ _03740_ _03616_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__or4b_1
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09448__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05788_ _01880_ _01881_ _01892_ net722 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a22o_2
XANTENNA__05470__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07161__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07527_ net450 _02840_ net442 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1078_X net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09463__A3 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07458_ core.register_file.registers_state\[831\] net683 _03562_ vssd1 vssd1 vccd1
+ vccd1 _03563_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06131__C1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08781__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05485__A1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06409_ net719 _02499_ _02507_ _02513_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__o22a_4
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07389_ net782 _03486_ _03492_ _03493_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_66_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09128_ _04805_ net2516 net350 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__mux2_1
XANTENNA__10632__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10230__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09059_ net611 _04855_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06985__B2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 core.register_file.registers_state\[262\] vssd1 vssd1 vccd1 vccd1 net1889
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 core.register_file.registers_state\[454\] vssd1 vssd1 vccd1 vccd1 net1900
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 core.ru.state\[6\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07529__A3 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__A1 core.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ clknet_leaf_4_clk _00533_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[493\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_109_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06737__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05645__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09687__A0 _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__A _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07162__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11854_ clknet_leaf_28_clk net50 net1194 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09439__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10805_ clknet_leaf_62_clk _00317_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[277\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11785_ clknet_leaf_28_clk _01289_ net1195 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08111__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07859__X _03964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10736_ clknet_leaf_106_clk _00248_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[208\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06899__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05476__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07578__Y _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ clknet_leaf_108_clk _00179_ net1135 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[139\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08414__A1 _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07217__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09611__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10598_ clknet_leaf_106_clk _00110_ net1158 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07100__A _03200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_131_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08178__B1 _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A1 core.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ clknet_leaf_97_clk _00731_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[691\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07754__B _03858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07076__S1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__07925__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__B2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09027__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05936__C1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06760_ core.register_file.registers_state\[529\] core.register_file.registers_state\[561\]
+ net883 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__mux2_1
XANTENNA__09678__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05951__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07770__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05711_ _01814_ _01815_ net618 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06691_ net805 _02794_ _02795_ net1084 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08585__B net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ net209 _04518_ net597 vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05642_ net1015 net898 _01507_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a21o_2
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08361_ _04453_ _04454_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05573_ net1042 core.register_file.registers_state\[859\] vssd1 vssd1 vccd1 vccd1
+ _01678_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07312_ _03416_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08292_ core.pc.current_pc\[6\] _04374_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06113__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07456__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09850__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload68_A clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07243_ _03346_ _03347_ net786 vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_95_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07174_ net995 core.register_file.registers_state\[579\] net883 core.register_file.registers_state\[611\]
+ net1079 vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07010__A _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06125_ net1051 core.register_file.registers_state\[456\] core.register_file.registers_state\[488\]
+ net677 net1015 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1038_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__A _02146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06056_ core.register_file.registers_state\[554\] core.register_file.registers_state\[522\]
+ net667 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout498_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 _05065_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_4
XANTENNA__08708__A2 _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout313 _05058_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06719__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
Xfanout335 _05046_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06719__B2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 _05027_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_2
XANTENNA__05465__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ net225 net2177 net380 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__mux2_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_4
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10090__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 _04898_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_4
XFILLER_0_94_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout379 net382 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_6
XANTENNA_fanout665_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ _04704_ net2030 net258 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__mux2_1
X_06958_ core.register_file.registers_state\[874\] core.register_file.registers_state\[842\]
+ net832 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
XANTENNA__09669__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__B2 core.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05909_ _02006_ _02007_ _02013_ _02010_ net964 net934 vssd1 vssd1 vccd1 vccd1 _02014_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09677_ _04876_ net292 net283 net2216 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout832_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06889_ net769 _02980_ _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__o21a_4
XANTENNA__10310__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ core.IO_mod.input_reg\[0\] net730 net249 _04691_ _04700_ vssd1 vssd1 vccd1
+ vccd1 _04703_ sky130_fd_sc_hd__o311ai_4
XANTENNA__06352__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08892__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ _04620_ _04622_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11570_ clknet_leaf_24_clk _01082_ net1187 vssd1 vssd1 vccd1 vccd1 core.decoder.inst\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09841__A0 _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ clknet_leaf_35_clk _00033_ net1220 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08942__C net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10452_ net1387 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07558__C _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06407__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10383_ net1406 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06502__S0 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09546__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08303__X _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input59_A gpio_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05630__B2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ clknet_leaf_43_clk _00516_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[476\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08175__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09372__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 net881 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__buf_2
Xfanout891 net894 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_4
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06591__C1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__A _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07135__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06343__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05697__A1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11837_ clknet_leaf_29_clk net63 net1199 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07589__X _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11768_ clknet_leaf_23_clk _01272_ net1187 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09832__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05449__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07989__A3 _04017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10719_ clknet_leaf_94_clk _00231_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11699_ clknet_leaf_76_clk _01211_ net1261 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06110__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06949__A1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07930_ _03922_ _03980_ _04034_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09899__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05285__A core.decoder.inst\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ _03414_ _03965_ _03418_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09600_ _04704_ net2432 net393 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06812_ net1066 _02911_ _02916_ net775 vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_88_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07792_ _03790_ _03869_ net477 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08596__A _03916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ _04877_ net399 net310 net2234 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a22o_1
X_06743_ _02816_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__or2_1
XANTENNA__07126__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09462_ _04958_ net320 net312 net2230 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06674_ net551 vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__inv_2
XANTENNA__07221__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08413_ core.pc.current_pc\[17\] _04498_ net229 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__o21ai_1
XANTENNA__05688__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06885__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05625_ _01722_ _01729_ net1026 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__mux2_1
X_09393_ net2206 net327 net316 _04861_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout246_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08344_ core.pc.current_pc\[11\] _04427_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05556_ net922 _01657_ _01658_ _01660_ net959 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__a311o_1
XFILLER_0_117_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08275_ core.pc.current_pc\[5\] _03231_ net577 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06101__A2 _02204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05487_ core.register_file.registers_state\[220\] core.register_file.registers_state\[252\]
+ net699 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout413_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07226_ core.register_file.registers_state\[545\] core.register_file.registers_state\[513\]
+ net849 vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07157_ net531 net504 _02518_ _01632_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06108_ net641 _02209_ _02210_ _02211_ _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07601__A2 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ net805 _03189_ _03188_ net790 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout782_A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05612__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06039_ net631 _02143_ net721 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a21o_1
XANTENNA__10305__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1110 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1110_X net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1208_X net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_4
XANTENNA__08157__A3 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07365__A1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07460__S1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05915__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09106__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _04930_ net289 net275 net2351 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07117__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10121__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06876__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10970__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__B net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ clknet_leaf_71_clk _01134_ net1270 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09814__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ clknet_leaf_27_clk _01065_ net1197 vssd1 vssd1 vccd1 vccd1 core.control_logic.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07569__B _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08093__A2 _04060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09290__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06723__S0 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ clknet_leaf_45_clk _00016_ net1288 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11326__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ clknet_leaf_41_clk _00996_ net1281 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[956\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10435_ net1449 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10188__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09276__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09593__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10366_ _05118_ net1621 net234 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05603__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10297_ net20 net905 _05244_ core.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 _01294_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09345__A2 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__A1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10360__A0 _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06564__C1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07108__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09024__B net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05410_ net924 net761 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08355__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06390_ net944 core.register_file.registers_state\[705\] net702 core.register_file.registers_state\[737\]
+ net643 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09805__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09040__A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05341_ wb.curr_state\[2\] wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__or2_4
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09281__A1 _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06095__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08060_ _02316_ _03201_ _03618_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05272_ net1123 core.control_logic.instruction\[5\] core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__and3b_1
XFILLER_0_114_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05842__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07011_ core.register_file.registers_state\[8\] core.register_file.registers_state\[40\]
+ core.register_file.registers_state\[136\] core.register_file.registers_state\[168\]
+ net872 net821 vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05842__B2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10179__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09584__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ _04849_ net738 vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__and2_1
X_07913_ net511 _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__nor2_2
X_08893_ net225 net737 vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__and2_1
X_07844_ net496 _03888_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10351__A0 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ _03787_ _03802_ net493 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__mux2_1
XANTENNA__07661__C _03231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10993__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ _04787_ net395 net307 net1874 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__a22o_1
X_06726_ net977 _02829_ _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06858__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09445_ _04924_ net315 net311 net2000 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a22o_1
X_06657_ core.register_file.registers_state\[852\] core.register_file.registers_state\[884\]
+ net888 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout530_A _03624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout628_A _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1272_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__B _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11349__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05608_ net1039 net748 core.register_file.registers_state\[791\] vssd1 vssd1 vccd1
+ vccd1 _01713_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09376_ net1865 net327 net315 _04770_ vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__a22o_1
X_06588_ net1106 core.register_file.registers_state\[726\] core.register_file.registers_state\[758\]
+ net852 net825 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08327_ _04421_ _04422_ _04419_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__o21a_1
X_05539_ net1034 core.register_file.registers_state\[474\] core.register_file.registers_state\[506\]
+ net670 net1010 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__o221a_1
XANTENNA__08075__A2 _03858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1060_X net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ core.pc.current_pc\[2\] core.pc.current_pc\[3\] vssd1 vssd1 vccd1 vccd1 _04362_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07209_ net994 core.register_file.registers_state\[322\] net884 core.register_file.registers_state\[354\]
+ net1078 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a221o_1
XANTENNA__05833__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ _01926_ _02840_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ net1127 net1442 net912 _05218_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__a31o_1
XANTENNA__05477__X _01582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05918__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09575__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ core.pc.current_pc\[30\] _05187_ _01386_ vssd1 vssd1 vccd1 vccd1 _05199_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09824__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ _04096_ net592 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07338__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07338__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08948__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10342__A0 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06546__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08667__C net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05910__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ clknet_leaf_13_clk _00496_ net1172 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[456\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09779__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06484__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11605_ clknet_leaf_27_clk _01117_ net1204 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10716__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08066__A2 _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09263__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07867__X _03972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09802__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07274__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ clknet_leaf_103_clk _01048_ net1156 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1008\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11467_ clknet_leaf_109_clk _00979_ net1134 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[939\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10866__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10418_ net1374 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08204__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11398_ clknet_leaf_99_clk _00910_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[870\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07577__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09019__B net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10349_ _05101_ net1811 net232 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
XANTENNA__05588__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09318__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07329__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07329__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09869__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10333__A0 _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05890_ _01991_ _01994_ net633 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06537__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06659__A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06001__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06001__B2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06511_ net973 _02614_ _02615_ net779 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__o31a_1
X_07491_ net1104 core.register_file.registers_state\[95\] core.register_file.registers_state\[127\]
+ net850 net810 vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07501__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09230_ _04807_ net421 net341 net1719 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06442_ core.register_file.registers_state\[153\] core.register_file.registers_state\[185\]
+ net714 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09161_ _04930_ net353 net343 net2194 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06373_ net647 _02476_ _02477_ net1031 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08112_ _03383_ _03384_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05324_ core.i_hit _01437_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__and2b_1
XANTENNA__07265__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ net2293 net365 net357 _04791_ vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05815__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08043_ _04059_ _04147_ net495 vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__mux2_1
XANTENNA__05815__B2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05255_ net1073 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold900 core.register_file.registers_state\[226\] vssd1 vssd1 vccd1 vccd1 net2219
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold911 core.register_file.registers_state\[510\] vssd1 vssd1 vccd1 vccd1 net2230
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout209_A _04334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05297__X _01412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold922 core.register_file.registers_state\[505\] vssd1 vssd1 vccd1 vccd1 net2241
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold933 core.pc.current_pc\[0\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08114__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold944 core.register_file.registers_state\[765\] vssd1 vssd1 vccd1 vccd1 net2263
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold955 core.register_file.registers_state\[690\] vssd1 vssd1 vccd1 vccd1 net2274
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 core.register_file.registers_state\[186\] vssd1 vssd1 vccd1 vccd1 net2285
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 core.register_file.registers_state\[126\] vssd1 vssd1 vccd1 vccd1 net2296
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1020_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 core.register_file.registers_state\[346\] vssd1 vssd1 vccd1 vccd1 net2307
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net1507 net541 net520 _02272_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__a22o_1
Xhold999 core.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06776__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1118_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06240__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08945_ net564 net215 net735 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout480_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout578_A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10324__A0 _05109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ net741 _04855_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_51_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ _03671_ _03674_ net505 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07758_ _03510_ _03812_ _03544_ _03480_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__o211a_1
XANTENNA__08784__A core.IO_mod.input_reg\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06709_ net550 _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout912_A _01449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ _01488_ _01550_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ net2199 net203 net405 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06700__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09359_ _05014_ net418 net412 net1712 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08048__A2 _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09245__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08008__B _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06059__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10889__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09819__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09796__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05806__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11321_ clknet_leaf_68_clk _00833_ net1267 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[793\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07847__B _02660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07008__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ clknet_leaf_57_clk _00764_ net1295 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[724\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07103__S0 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ net93 net919 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08756__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ clknet_leaf_83_clk _00695_ net1231 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[655\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08959__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09554__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A gpio_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _05183_ _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05665__S0 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08678__B _04746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10065_ _04186_ net592 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__nand2_1
XANTENNA__10315__A0 _05100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06519__C1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09720__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__C1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06090__S0 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10967_ clknet_leaf_20_clk _00479_ net1188 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[439\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10898_ clknet_leaf_69_clk _00410_ net1277 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[370\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09787__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11519_ clknet_leaf_41_clk _01031_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[991\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold207 _01223_ vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 core.register_file.registers_state\[403\] vssd1 vssd1 vccd1 vccd1 net1537
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 core.IO_mod.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06470__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05558__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06470__B2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout709 net711 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08869__A _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06991_ net1100 core.register_file.registers_state\[329\] core.register_file.registers_state\[361\]
+ net844 net980 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__o221a_1
XANTENNA__07970__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05430__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08588__B net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ net608 net220 vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__and2_2
XANTENNA__10306__A0 _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05942_ net945 core.register_file.registers_state\[334\] net705 core.register_file.registers_state\[366\]
+ net1017 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09172__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1280 net1281 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__clkbuf_4
Xfanout1291 net1292 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__clkbuf_4
X_08661_ net1979 net469 net438 _04732_ vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__a22o_1
X_05873_ net629 _01968_ _01971_ _01966_ net718 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__o311a_2
X_07612_ _03714_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__nand2_1
X_08592_ _01435_ net474 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_89_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05733__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07543_ net507 _03645_ _03647_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_49_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08598__D_N _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06289__A1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09212__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ net1028 _03575_ _03578_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08683__C1 _04750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05497__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09213_ net571 _04707_ net422 net342 net1721 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__a32o_1
X_06425_ _02527_ _02528_ _01895_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__or3b_4
XFILLER_0_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09227__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09144_ _04714_ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout1068_A core.decoder.inst\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06356_ net952 core.register_file.registers_state\[66\] net710 core.register_file.registers_state\[98\]
+ net661 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a221o_1
XANTENNA__08543__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05307_ core.d_hit net731 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09075_ net1121 net606 vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06287_ _02389_ _02391_ net619 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06997__C1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold730 core.register_file.registers_state\[496\] vssd1 vssd1 vccd1 vccd1 net2049
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold741 core.register_file.registers_state\[44\] vssd1 vssd1 vccd1 vccd1 net2060
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout695_A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 core.register_file.registers_state\[504\] vssd1 vssd1 vccd1 vccd1 net2071
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold763 core.register_file.registers_state\[236\] vssd1 vssd1 vccd1 vccd1 net2082
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 core.register_file.registers_state\[433\] vssd1 vssd1 vccd1 vccd1 net2093
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1023_X net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 core.register_file.registers_state\[251\] vssd1 vssd1 vccd1 vccd1 net2104
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11537__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 core.register_file.registers_state\[254\] vssd1 vssd1 vccd1 vccd1 net2115
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09977_ net1129 net1632 net893 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout862_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net2126 net367 _04925_ net431 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__a22o_1
XANTENNA__06299__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07970__X _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09163__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ _04780_ net2371 net372 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07174__C1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06072__S0 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ clknet_leaf_53_clk _01339_ net1300 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11136__RESET_B net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10821_ clknet_leaf_87_clk _00333_ net1229 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[293\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08945__C net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10076__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10752_ clknet_leaf_51_clk _00264_ net1304 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[224\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08019__A _03397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10268__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ clknet_leaf_25_clk _00195_ net1186 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[155\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07229__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09549__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__A2 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05378__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ clknet_leaf_13_clk _00816_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[776\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08729__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11235_ clknet_leaf_64_clk _00747_ net1248 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[707\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09284__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10000__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ clknet_leaf_95_clk _00678_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[638\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05412__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ _03884_ _03945_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__nor2_1
X_11097_ clknet_leaf_68_clk _00609_ net1265 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[569\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05963__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__X _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10048_ _05123_ net515 vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__nor2_4
XANTENNA__06002__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07165__C1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold90 core.register_file.registers_state\[967\] vssd1 vssd1 vccd1 vccd1 net1409
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07704__B2 _03808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08901__B1 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06063__S0 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05715__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10067__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10859__RESET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08680__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06210_ net554 _02314_ _02278_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07768__A _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07190_ net995 core.register_file.registers_state\[962\] net883 core.register_file.registers_state\[994\]
+ net983 vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06141_ core.register_file.registers_state\[7\] net705 net644 _02245_ vssd1 vssd1
+ vccd1 vccd1 _02246_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06072_ core.register_file.registers_state\[777\] core.register_file.registers_state\[809\]
+ core.register_file.registers_state\[905\] core.register_file.registers_state\[937\]
+ net701 net1015 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09900_ _05004_ net388 net377 net2286 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08196__A1 _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout506 net509 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_2
XANTENNA__09393__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout517 _05126_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08735__A3 _04794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ net216 net2053 net381 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
Xfanout528 _03625_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_8
Xfanout539 _01631_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10584__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ _04993_ net289 net257 net1775 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__a22o_1
X_06974_ net775 _03072_ _03073_ net771 vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a31o_1
XANTENNA__05954__B1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08713_ net563 net431 _04776_ net466 net1577 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__a32o_1
X_05925_ net927 _02029_ _02028_ net1006 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_33_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _04890_ net2217 net278 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
XANTENNA__08499__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ _01620_ _04662_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__or2_2
XFILLER_0_96_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05856_ core.register_file.registers_state\[17\] net689 net661 _01960_ vssd1 vssd1
+ vccd1 vccd1 _01961_ sky130_fd_sc_hd__a211o_1
XANTENNA__05706__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05751__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08575_ _01418_ _01618_ _01629_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05787_ _01886_ _01891_ _01521_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout443_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07526_ net454 net446 vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06285__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07457_ core.register_file.registers_state\[799\] net700 vssd1 vssd1 vccd1 vccd1
+ _03562_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout610_A _04669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__A2 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08781__B net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout708_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ net633 _02509_ _02512_ net723 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07388_ net788 _03488_ _03489_ net782 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a31o_1
X_09127_ net218 net2280 net347 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__mux2_1
X_06339_ _02440_ _02443_ net630 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__o21a_1
XANTENNA__10308__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09058_ net1001 net464 _05011_ net430 net1946 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08009_ _02206_ _03111_ net579 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold560 core.register_file.registers_state\[820\] vssd1 vssd1 vccd1 vccd1 net1879
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 net160 vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ clknet_leaf_101_clk _00532_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[492\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold582 core.register_file.registers_state\[632\] vssd1 vssd1 vccd1 vccd1 net1901
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold593 core.register_file.registers_state\[788\] vssd1 vssd1 vccd1 vccd1 net1912
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05945__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__A0 _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09832__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07352__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11853_ clknet_leaf_36_clk net49 net1221 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06370__B1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ clknet_leaf_55_clk _00316_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[276\]
+ sky130_fd_sc_hd__dfrtp_1
X_11784_ clknet_leaf_29_clk _01288_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08972__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ clknet_leaf_82_clk _00247_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[207\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_40_clk_X clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__A2 _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09279__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06673__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08618__C_N _03964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ clknet_leaf_106_clk _00178_ net1138 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[138\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11702__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10597_ clknet_leaf_87_clk _00109_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_55_clk_X clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05395__X _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ clknet_leaf_67_clk _00730_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[690\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09375__B1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06431__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06189__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__07386__C1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
X_11149_ clknet_leaf_4_clk _00661_ net1141 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[621\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09027__B net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05936__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05710_ net948 core.register_file.registers_state\[149\] net763 net928 vssd1 vssd1
+ vccd1 vccd1 _01815_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06690_ net988 core.register_file.registers_state\[691\] net869 core.register_file.registers_state\[659\]
+ net817 vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__o221a_1
XANTENNA__09043__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05641_ net555 _01745_ _01711_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08360_ _04431_ _04435_ _04445_ _04453_ _04443_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__o311a_1
XANTENNA__05290__B _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05572_ net937 core.register_file.registers_state\[891\] net758 vssd1 vssd1 vccd1
+ vccd1 _01677_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10693__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07311_ _02751_ _02783_ _02750_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_138_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08291_ _04378_ _04388_ _04389_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_138_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09850__A1 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06664__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ net990 core.register_file.registers_state\[65\] net876 core.register_file.registers_state\[97\]
+ net824 vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a221o_1
XANTENNA__06664__B2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05872__C1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07173_ core.register_file.registers_state\[547\] core.register_file.registers_state\[515\]
+ net855 vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07785__X _03890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09917__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06124_ net1051 core.register_file.registers_state\[328\] core.register_file.registers_state\[360\]
+ net677 net925 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07613__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06055_ _02156_ _02159_ net717 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07945__B _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09366__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 net306 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_6
XFILLER_0_26_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09905__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout314 _05058_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_4
XANTENNA__07916__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout393_A _05066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout336 _05046_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_4
Xfanout347 _05025_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_6
X_09814_ net226 net2416 net381 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
Xfanout358 net362 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_4
XANTENNA__09118__A0 _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 _04898_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_6
XFILLER_0_96_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _04961_ net290 vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__nand2_1
X_06957_ core.register_file.registers_state\[810\] core.register_file.registers_state\[778\]
+ net832 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout560_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05908_ _02011_ _02012_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__and2_1
X_06888_ net777 _02987_ _02992_ net773 vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09676_ _04871_ net290 net283 net2379 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__a22o_1
X_08627_ _01621_ _03739_ _04698_ _04699_ _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__o221ai_4
X_05839_ core.register_file.registers_state\[16\] core.register_file.registers_state\[48\]
+ net695 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06352__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08558_ _04633_ _04634_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07509_ _03612_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__xnor2_1
X_08489_ net1124 _03536_ net574 vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10520_ clknet_leaf_35_clk _00032_ net1220 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10451_ net1340 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09827__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ net1470 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06502__S1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11105__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold390 core.register_file.registers_state\[568\] vssd1 vssd1 vccd1 vccd1 net1709
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ clknet_leaf_25_clk _00515_ net1191 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[475\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09562__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06186__A3 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
XANTENNA__09109__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_4
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11255__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07590__B _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06487__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07082__S _01462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1090 core.register_file.registers_state\[223\] vssd1 vssd1 vccd1 vccd1 net2409
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06343__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11836_ clknet_leaf_29_clk net62 net1195 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06493__Y _02598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ clknet_leaf_28_clk _01271_ net1194 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05449__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ clknet_leaf_96_clk _00230_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[190\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11698_ clknet_leaf_49_clk net1524 net1309 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05854__C1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_20_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ clknet_leaf_54_clk _00161_ net1298 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09596__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__A _02146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06949__A2 _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07257__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09348__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _03413_ _03416_ _03419_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05853__X _01958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06811_ _02912_ _02913_ _02914_ _02915_ net978 net1083 vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__mux4_1
X_07791_ net488 _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06582__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06742_ _02845_ _02846_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09530_ _04872_ net457 net307 net2045 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09520__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _04956_ net316 net311 net2051 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a22o_1
X_06673_ net769 _02777_ _02765_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06334__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05732__C net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ core.pc.current_pc\[17\] _04498_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__and2_2
XANTENNA__06885__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05624_ net933 _01723_ _01724_ _01727_ _01728_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__o32a_1
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09392_ net1701 net327 net316 _04856_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08343_ core.pc.current_pc\[10\] _04439_ net597 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08087__B1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05555_ net938 core.register_file.registers_state\[1018\] net757 _01659_ net1010
+ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__o311a_1
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_108_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout239_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06098__C1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06637__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _04366_ _04368_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06637__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05486_ core.register_file.registers_state\[156\] core.register_file.registers_state\[188\]
+ net699 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07225_ net1086 _03326_ _03329_ net1068 vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__o211ai_1
XANTENNA__07021__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1050_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__A _03826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06107_ net942 core.register_file.registers_state\[680\] net751 net1013 vssd1 vssd1
+ vccd1 vccd1 _02212_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_37_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07062__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07087_ _03190_ _03191_ net784 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a21o_1
XANTENNA__07062__B2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1315_A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09339__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06038_ net958 _02137_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout775_A _01463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1103_X net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05376__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout942_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ net511 _03957_ _04017_ _04091_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05376__B2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _04928_ net295 net276 net1895 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05415__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09511__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _04781_ net289 net283 net2211 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__a22o_1
XANTENNA__08793__Y _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__RESET_B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06876__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07630__S net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11621_ clknet_leaf_76_clk _01133_ net1260 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06628__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ clknet_leaf_33_clk _01064_ net1208 vssd1 vssd1 vccd1 vccd1 core.control_logic.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07569__C net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06723__S1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10503_ clknet_leaf_46_clk _00015_ net1290 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11483_ clknet_leaf_22_clk _00995_ net1181 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[955\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09578__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ net1394 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09557__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06770__A _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07053__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10365_ _05117_ net1506 net235 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07077__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05603__A2 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10296_ net19 net902 net796 net1678 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07805__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05367__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05367__B2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08305__A1 _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10112__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10795__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05552__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11819_ clknet_leaf_48_clk _01320_ net1312 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09805__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05340_ wb.curr_state\[2\] wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09040__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05827__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05271_ core.pc.current_pc\[31\] vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07010_ _03111_ _03114_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__nor2_1
XANTENNA__09569__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11420__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08792__A1 core.IO_mod.input_reg\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08961_ net2308 net367 _04947_ net431 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ _02385_ _03684_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__or2_4
X_08892_ net2506 net369 _04901_ net436 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__a22o_1
XANTENNA__05583__X _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09741__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ net491 _03906_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07774_ _03750_ _03782_ net494 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__mux2_2
XANTENNA__08894__X _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09513_ _04782_ net397 net308 net1956 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__a22o_1
X_06725_ net1110 core.register_file.registers_state\[978\] core.register_file.registers_state\[1010\]
+ net851 net1080 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o221a_1
XANTENNA__10103__A1 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout356_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _04922_ net318 net311 net1846 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__a22o_1
X_06656_ core.register_file.registers_state\[788\] core.register_file.registers_state\[820\]
+ net888 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07450__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05607_ net1039 net748 core.register_file.registers_state\[919\] vssd1 vssd1 vccd1
+ vccd1 _01712_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_23_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06587_ net1106 core.register_file.registers_state\[598\] core.register_file.registers_state\[630\]
+ net852 net810 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_23_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09375_ net1986 net327 net319 _04764_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1265_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08326_ _04419_ _04421_ _04422_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nor3_1
X_05538_ net1034 core.register_file.registers_state\[346\] core.register_file.registers_state\[378\]
+ net670 net922 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10518__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ core.pc.current_pc\[2\] core.pc.current_pc\[3\] vssd1 vssd1 vccd1 vccd1 _04361_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05469_ net1051 core.register_file.registers_state\[221\] core.register_file.registers_state\[253\]
+ net677 net664 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07208_ core.register_file.registers_state\[290\] core.register_file.registers_state\[258\]
+ core.register_file.registers_state\[418\] core.register_file.registers_state\[386\]
+ net856 net1078 vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__mux4_1
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08188_ net546 _04292_ net901 _01896_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout892_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07139_ net994 core.register_file.registers_state\[324\] net884 core.register_file.registers_state\[356\]
+ net1078 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10316__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08783__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ core.pc.current_pc\[30\] _01386_ _05187_ vssd1 vssd1 vccd1 vccd1 _05198_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_112_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__C1 _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07692__Y _03797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ core.pc.current_pc\[12\] net590 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__or2_1
XANTENNA__07625__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08948__C net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06101__Y _02206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09840__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10983_ clknet_leaf_93_clk _00495_ net1237 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08838__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11604_ clknet_leaf_29_clk _01116_ net1198 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09799__B1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08980__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07274__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11535_ clknet_leaf_79_clk _01047_ net1251 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1007\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09287__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07596__A _02530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06482__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11466_ clknet_leaf_1_clk _00978_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[938\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07026__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10417_ net1341 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07026__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11397_ clknet_leaf_86_clk _00909_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08204__B _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10030__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05588__A1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10348_ _05100_ net1563 net233 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__mux2_1
XANTENNA__09019__C net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ net32 net904 net797 core.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__a22o_1
XANTENNA__08526__A1 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09723__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10097__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06510_ net1096 core.register_file.registers_state\[349\] core.register_file.registers_state\[381\]
+ net838 net981 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_66_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07490_ core.register_file.registers_state\[31\] core.register_file.registers_state\[63\]
+ core.register_file.registers_state\[159\] core.register_file.registers_state\[191\]
+ net873 net822 vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__mux4_1
XANTENNA__06675__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07270__S net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06441_ _02540_ _02545_ net634 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__mux2_1
XANTENNA__09051__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ _04928_ net358 net345 net2170 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09986__A _05096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06372_ core.register_file.registers_state\[674\] net688 net661 _02474_ vssd1 vssd1
+ vccd1 vccd1 _02477_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08890__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09254__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ _03383_ _03384_ net530 vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05323_ _01429_ _01432_ _01436_ net34 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__o31a_1
XANTENNA__07265__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ net2176 net363 net351 _04786_ vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__a22o_1
XANTENNA__06699__S0 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08042_ net486 _04117_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05254_ net1111 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XANTENNA__06473__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05371__S0 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold901 core.register_file.registers_state\[460\] vssd1 vssd1 vccd1 vccd1 net2220
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 core.register_file.registers_state\[155\] vssd1 vssd1 vccd1 vccd1 net2231
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07017__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07017__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold923 core.register_file.registers_state\[631\] vssd1 vssd1 vccd1 vccd1 net2242
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold934 core.register_file.registers_state\[449\] vssd1 vssd1 vccd1 vccd1 net2253
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 core.register_file.registers_state\[462\] vssd1 vssd1 vccd1 vccd1 net2264
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07656__D net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08765__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__X _03898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06225__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 core.register_file.registers_state\[216\] vssd1 vssd1 vccd1 vccd1 net2275
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold967 core.register_file.registers_state\[917\] vssd1 vssd1 vccd1 vccd1 net2286
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 core.register_file.registers_state\[923\] vssd1 vssd1 vccd1 vccd1 net2297
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net1581 net540 net519 _02314_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__a22o_1
Xhold989 core.register_file.registers_state\[120\] vssd1 vssd1 vccd1 vccd1 net2308
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10960__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06240__A2 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08944_ _04815_ net735 vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_55_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1013_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09714__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ net211 net2450 net374 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout473_A _05127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07826_ net1112 _03928_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07757_ net529 _03841_ _03842_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout640_A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ _01895_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07688_ core.decoder.inst\[30\] net900 net546 _03792_ vssd1 vssd1 vccd1 vccd1 _03793_
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__06585__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09599__C net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A2 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07033__X _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09427_ net1915 net210 net407 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XANTENNA__05503__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06639_ net1087 _02740_ _02743_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05503__B2 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07968__X _04073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09358_ _05013_ net416 net412 net1783 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09245__A2 _04851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ _02207_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ net2192 _04895_ net335 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11320_ clknet_leaf_2_clk _00832_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[792\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06464__C1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ clknet_leaf_10_clk _00763_ net1149 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[723\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08799__X _04849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__RESET_B net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07103__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06216__C1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ net1128 net1627 net913 _05209_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a31o_1
XANTENNA__09835__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__B2 _04812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ clknet_leaf_81_clk _00694_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[654\]
+ sky130_fd_sc_hd__dfrtp_1
X_10133_ core.pc.current_pc\[28\] _05178_ net588 vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08959__B net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05665__S1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ core.pc.current_pc\[5\] net591 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__or2_1
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05990__A1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06519__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06090__S1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06495__A _02534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ clknet_leaf_60_clk _00478_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[438\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09484__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10897_ clknet_leaf_66_clk _00409_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[369\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09236__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ clknet_leaf_94_clk _01030_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[990\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06434__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08215__A _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold208 core.register_file.registers_state\[915\] vssd1 vssd1 vccd1 vccd1 net1527
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 net171 vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10983__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11449_ clknet_leaf_64_clk _00961_ net1249 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[921\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08747__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06207__C1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08869__B _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06990_ net1100 core.register_file.registers_state\[457\] core.register_file.registers_state\[489\]
+ net843 net1074 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11339__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05574__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05430__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09046__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05941_ net1029 _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__or2_1
XANTENNA__05981__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05981__B2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1270 net1271 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_68_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05872_ net660 _01975_ _01976_ net618 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__o211a_1
X_08660_ net572 net609 net224 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__and3_1
Xfanout1281 net1283 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_2
Xfanout1292 net1313 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__buf_2
XANTENNA__08885__A core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__A2 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ net454 _03289_ net446 net498 vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08591_ _01504_ _04651_ _04665_ _01422_ net34 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__o2111a_4
XANTENNA__05733__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07542_ net502 _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09475__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ net961 _03576_ _03577_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__or3_1
XANTENNA__07486__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ net1121 net605 _05030_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__or3_4
X_06424_ _02527_ _02528_ _01895_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_8_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09227__A2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06355_ _02457_ _02459_ net619 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_44_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ net1121 net735 vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05306_ core.d_hit net727 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06446__C1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09074_ net998 net463 _05021_ net428 net1795 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__a32o_1
X_06286_ core.register_file.registers_state\[3\] net710 net647 _02390_ vssd1 vssd1
+ vccd1 vccd1 _02391_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08025_ _04080_ _04088_ net487 vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1130_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold720 core.register_file.registers_state\[356\] vssd1 vssd1 vccd1 vccd1 net2039
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 core.register_file.registers_state\[381\] vssd1 vssd1 vccd1 vccd1 net2050
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09935__A0 core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold742 core.register_file.registers_state\[214\] vssd1 vssd1 vccd1 vccd1 net2061
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1228_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold753 core.register_file.registers_state\[179\] vssd1 vssd1 vccd1 vccd1 net2072
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 core.register_file.registers_state\[580\] vssd1 vssd1 vccd1 vccd1 net2083
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08412__X _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold775 core.register_file.registers_state\[319\] vssd1 vssd1 vccd1 vccd1 net2094
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 core.register_file.registers_state\[107\] vssd1 vssd1 vccd1 vccd1 net2105
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold797 core.IO_mod.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09976_ core.d_hit _01367_ _01441_ _01445_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1016_X net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05421__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05484__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ net563 _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__and2_1
XANTENNA__05972__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05972__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ net222 core.register_file.registers_state\[75\] net371 vssd1 vssd1 vccd1
+ vccd1 _00115_ sky130_fd_sc_hd__mux2_1
XANTENNA__08795__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07174__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ net511 _03909_ _03913_ _03658_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a211o_1
XANTENNA__08910__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05724__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06072__S1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05724__B2 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08789_ net462 _04711_ _04840_ net466 net2444 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__a32o_1
X_10820_ clknet_leaf_77_clk _00332_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09466__A2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07477__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ clknet_leaf_94_clk _00263_ net1240 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[223\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11176__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06685__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09218__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10682_ clknet_leaf_7_clk _00194_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[154\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07229__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__A3 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06254__S net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08035__A _04139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11303_ clknet_leaf_91_clk _00815_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[775\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09926__A0 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09565__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ clknet_leaf_80_clk _00746_ net1253 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[706\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11165_ clknet_leaf_19_clk _00677_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[637\]
+ sky130_fd_sc_hd__dfrtp_1
X_10116_ net470 _05168_ _05169_ net515 net1436 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a32o_1
X_11096_ clknet_leaf_10_clk _00608_ net1149 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[568\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ _05122_ _05124_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_106_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold80 core.register_file.registers_state\[6\] vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07704__A2 _03788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold91 core.register_file.registers_state\[992\] vssd1 vssd1 vccd1 vccd1 net1410
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_102_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08901__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06063__S1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05715__A1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11781__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09457__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10949_ clknet_leaf_100_clk _00461_ net1165 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[421\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05479__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09209__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11011__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07401__X _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__B _03476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06140_ net945 core.register_file.registers_state\[39\] net766 vssd1 vssd1 vccd1
+ vccd1 _02245_ sky130_fd_sc_hd__or3_1
XANTENNA__10899__RESET_B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09090__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06071_ net583 _02174_ _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_77_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09917__A0 core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05651__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10729__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout507 net509 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_4
X_09830_ net217 net1975 net380 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
Xfanout518 _05126_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_2
Xfanout529 _03624_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_4
XANTENNA__05403__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06600__C1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ _04991_ net294 net258 net1888 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05735__C net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06973_ net1083 _03074_ _03077_ net779 vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__o211a_1
XANTENNA__08886__Y _04897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__A1 _04705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ net606 net222 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2_2
X_05924_ net947 core.register_file.registers_state\[974\] net705 core.register_file.registers_state\[1006\]
+ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09692_ net206 net1909 net279 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10879__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08643_ _01620_ _04662_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nor2_2
X_05855_ net1059 core.register_file.registers_state\[49\] net755 vssd1 vssd1 vccd1
+ vccd1 _01960_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08574_ core.pc.current_pc\[31\] _04649_ net595 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09448__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05786_ net620 _01890_ _01889_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07525_ _01613_ _02525_ _03627_ _03628_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_46_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1080_A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout436_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1178_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06131__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ core.register_file.registers_state\[991\] net707 _03551_ vssd1 vssd1 vccd1
+ vccd1 _03561_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06131__B2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08781__C net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06407_ _02510_ _02511_ net963 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a21o_1
XANTENNA__05485__A3 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ _03490_ _03491_ net793 vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05890__B1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11504__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ net219 net2349 net349 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__mux2_1
X_06338_ net624 _02441_ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09081__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07965__Y _04070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06269_ net952 core.register_file.registers_state\[452\] vssd1 vssd1 vccd1 vccd1
+ _02374_ sky130_fd_sc_hd__and2_1
X_09057_ net744 net613 net211 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__and3_1
XANTENNA__10230__A3 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ _02206_ _03111_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__nand2_1
XANTENNA__05642__B1 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09908__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold550 core.register_file.registers_state\[572\] vssd1 vssd1 vccd1 vccd1 net1869
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 core.register_file.registers_state\[582\] vssd1 vssd1 vccd1 vccd1 net1880
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout972_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 core.register_file.registers_state\[491\] vssd1 vssd1 vccd1 vccd1 net1891
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 core.register_file.registers_state\[408\] vssd1 vssd1 vccd1 vccd1 net1902
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10324__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06198__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 core.register_file.registers_state\[436\] vssd1 vssd1 vccd1 vccd1 net1913
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08302__B _04401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06103__A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ net1451 net2554 net798 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05645__C net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07490__S0 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05945__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08895__B1 _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11852_ clknet_leaf_37_clk net48 net1223 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09439__A2 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ clknet_leaf_98_clk _00315_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[275\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08647__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11783_ clknet_leaf_24_clk _01287_ net1183 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08972__B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10734_ clknet_leaf_89_clk _00246_ net1233 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[206\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10665_ clknet_leaf_40_clk _00177_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[137\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ clknet_leaf_76_clk _00108_ net1260 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09611__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07083__C1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05676__X _01781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05633__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08178__A2 _03949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11217_ clknet_leaf_74_clk _00729_ net1257 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[689\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06189__A1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_78_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11148_ clknet_leaf_103_clk _00660_ net1156 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[620\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05936__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ clknet_leaf_90_clk _00591_ net1243 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[551\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09678__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07233__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09043__B net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05640_ net721 _01730_ _01738_ _01744_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__o2bb2a_4
XTAP_TAPCELL_ROW_86_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11027__RESET_B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05571_ net1004 _01672_ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07310_ _02691_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__nand2_1
XANTENNA__06649__C1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11527__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08290_ net230 _04390_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__nor2_1
XANTENNA__06683__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09850__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07241_ net991 core.register_file.registers_state\[193\] net877 core.register_file.registers_state\[225\]
+ net808 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a221o_1
XANTENNA__05299__A core.decoder.inst\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07172_ net995 core.register_file.registers_state\[643\] net883 core.register_file.registers_state\[675\]
+ net983 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06123_ core.register_file.registers_state\[264\] core.register_file.registers_state\[296\]
+ core.register_file.registers_state\[392\] core.register_file.registers_state\[424\]
+ net701 net1015 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux4_1
XANTENNA__10551__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07613__A1 _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__A3 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06054_ net1025 _02157_ _02158_ net628 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a31o_1
XANTENNA__06821__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06622__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08169__A2 _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09366__B2 _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08122__B _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08897__X _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout315 net317 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout326 _05056_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_4
X_09813_ net207 net2387 net380 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07019__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout337 _05046_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_6
XFILLER_0_96_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout348 _05025_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_4
XANTENNA__05465__C net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout359 net361 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_4
XANTENNA_fanout386_A _05085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net241 net736 net290 net275 net1829 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__a32o_1
X_06956_ _03057_ _03058_ _03060_ _03059_ net789 net802 vssd1 vssd1 vccd1 vccd1 _03061_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09669__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05907_ net951 core.register_file.registers_state\[719\] net709 core.register_file.registers_state\[751\]
+ net646 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a221o_1
X_09675_ _04866_ net292 net284 net2315 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__a22o_1
X_06887_ net1087 _02988_ _02991_ net783 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout1295_A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _04700_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__inv_2
XANTENNA__06888__C1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05838_ net1037 core.register_file.registers_state\[176\] net668 core.register_file.registers_state\[144\]
+ net637 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a221o_1
XANTENNA__06352__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ _01488_ _04335_ _04630_ _01508_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05769_ net617 _01872_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_X net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07689__A _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07508_ _01550_ _02602_ _01632_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08284__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08488_ core.pc.current_pc\[23\] net600 _04570_ _04571_ vssd1 vssd1 vccd1 vccd1 _00031_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08137__X _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07439_ _03509_ _03542_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nand2_1
XANTENNA__10319__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1250_X net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10450_ net1388 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07065__C1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ net607 net242 net356 net364 net1752 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__a32o_1
X_10381_ net1446 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05615__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout975_X net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09357__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 core.register_file.registers_state\[786\] vssd1 vssd1 vccd1 vccd1 net1699
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 core.register_file.registers_state\[429\] vssd1 vssd1 vccd1 vccd1 net1710
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09843__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ clknet_leaf_6_clk _00514_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[474\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09109__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
Xfanout871 net874 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_4
Xfanout882 _01457_ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_2
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06591__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__A0 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1080 core.register_file.registers_state\[206\] vssd1 vssd1 vccd1 vccd1 net2399
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_88_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1091 core.register_file.registers_state\[99\] vssd1 vssd1 vccd1 vccd1 net2410
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08983__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__X _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11835_ clknet_leaf_36_clk net61 net1221 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11766_ clknet_leaf_28_clk _01270_ net1194 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09293__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10717_ clknet_leaf_17_clk _00229_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[189\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ clknet_leaf_72_clk net1477 net1269 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05854__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10648_ clknet_leaf_3_clk _00160_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10579_ clknet_leaf_96_clk _00091_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06442__S net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05701__S0 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09348__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06031__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06810_ net1092 core.register_file.registers_state\[845\] core.register_file.registers_state\[877\]
+ net831 vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__o22a_1
XANTENNA__08369__S net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ net477 _03892_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_88_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07126__X _03231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09054__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06741_ _02840_ _02844_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nand2_1
XANTENNA__08859__A0 _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09520__A1 _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ _04954_ net322 net313 net1981 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__a22o_1
X_06672_ net781 _02770_ _02771_ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__o31a_1
XANTENNA__08893__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08411_ core.pc.current_pc\[16\] net598 _04501_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05623_ net638 _01725_ _01726_ net1004 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a31o_1
XANTENNA__05688__A3 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09391_ net1853 net329 net324 _04850_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08342_ _04438_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__inv_2
XANTENNA__08087__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05554_ net1039 core.register_file.registers_state\[986\] vssd1 vssd1 vccd1 vccd1
+ _01659_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08273_ core.pc.current_pc\[5\] _04370_ net230 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09995__Y _05098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05485_ net950 core.register_file.registers_state\[380\] net764 _01589_ net927 vssd1
+ vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__o311a_1
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09928__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ _03327_ _03328_ net974 vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05940__S0 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07047__C1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__B _04018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _03247_ _03248_ _03259_ net770 vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__o22a_4
XANTENNA_fanout301_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06106_ net1046 net751 core.register_file.registers_state\[648\] vssd1 vssd1 vccd1
+ vccd1 _02211_ sky130_fd_sc_hd__a21o_1
XANTENNA__07448__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07086_ net988 core.register_file.registers_state\[198\] net871 core.register_file.registers_state\[230\]
+ net805 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a221o_1
X_06037_ _02138_ _02139_ _02141_ net923 net1025 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1210_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1308_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08011__B2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__B _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07988_ net1112 _04090_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _04926_ net295 net276 net1955 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__a22o_1
X_06939_ net1083 _03042_ _03043_ net968 vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _04776_ net288 net282 net1831 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07911__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ _04278_ _04306_ _04317_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _04943_ net401 net300 net2202 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11620_ clknet_leaf_49_clk _01132_ net1310 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07825__A1 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11551_ clknet_leaf_41_clk _01063_ net1279 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1023\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06184__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ clknet_leaf_46_clk _00014_ net1290 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[6\]
+ sky130_fd_sc_hd__dfrtp_2
Xwire524 _05097_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_2
XANTENNA__09838__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire535 _02380_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_4
X_11482_ clknet_leaf_7_clk _00994_ net1145 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[954\]
+ sky130_fd_sc_hd__dfstp_1
X_10433_ net1368 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10188__A2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__B1 _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A gpio_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ _05116_ net1682 net233 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__mux2_1
XANTENNA__05603__A3 _01706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10295_ net18 net904 net797 net2515 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__a22o_1
XANTENNA__08978__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07210__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06498__A _01550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06564__A1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout690 net691 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_2
XANTENNA__05772__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07821__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11818_ clknet_leaf_50_clk _01319_ net1307 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06437__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09805__A2 _04851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ clknet_leaf_32_clk _01261_ net1207 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09040__C net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05270_ core.pc.current_pc\[28\] vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XANTENNA__06095__A3 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09569__A1 _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__A2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09049__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06252__B1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ net563 net212 net735 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08888__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07911_ _04012_ _04015_ net490 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__mux2_2
XANTENNA__06900__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ net569 net226 net739 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__and3_1
XANTENNA__07201__C1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ _03449_ _03541_ _03545_ _03547_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or4_1
XANTENNA_wire524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ net265 _03872_ _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09512_ net564 _04776_ net395 net307 net1609 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__a32o_1
X_06724_ net1110 core.register_file.registers_state\[850\] core.register_file.registers_state\[882\]
+ net860 net984 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06307__A1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10103__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09443_ _04920_ net315 net311 net1891 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06655_ core.register_file.registers_state\[980\] core.register_file.registers_state\[1012\]
+ net888 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout349_A _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05606_ net583 _01710_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09374_ net1887 net328 net319 _04759_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__a22o_1
XANTENNA__09257__B1 _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06586_ net552 _02689_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08325_ _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05537_ net1025 _01641_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout516_A _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1160_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1258_A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05818__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ net231 net596 vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__and2b_4
XANTENNA__08480__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05468_ net1051 core.register_file.registers_state\[93\] core.register_file.registers_state\[125\]
+ net677 net641 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11245__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07207_ net792 _03310_ _03311_ _03309_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__a31o_1
XANTENNA__06491__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _01926_ _02840_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05399_ _01495_ _01503_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__RESET_B net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07178__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07138_ core.register_file.registers_state\[292\] core.register_file.registers_state\[260\]
+ core.register_file.registers_state\[420\] core.register_file.registers_state\[388\]
+ net856 net1078 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__mux4_1
XANTENNA__05918__C net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__A2 _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07069_ _02276_ _03173_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06794__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1213_X net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11395__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10080_ net472 _05146_ _05147_ net517 net1442 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__a32o_1
XANTENNA__08150__X _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__S net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06546__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ clknet_leaf_98_clk _00494_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[454\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09496__B1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05950__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06257__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09248__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ clknet_leaf_25_clk _01115_ net1193 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09799__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07259__C1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08980__B net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05809__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11534_ clknet_leaf_90_clk _01046_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1006\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ clknet_leaf_17_clk _00977_ net1211 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[937\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05397__A _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__C1 _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ net1324 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11396_ clknet_leaf_81_clk _00908_ net1255 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10030__B2 _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07577__A3 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10347_ _05099_ net1532 net234 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06785__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06785__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10278_ net31 net903 net795 net2522 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__o22a_1
XANTENNA__05993__C1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_107_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06537__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__B1 _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06537__B2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05745__C1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05563__C net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09487__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10097__A1 _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05860__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06440_ _02541_ _02542_ _02543_ _02544_ net648 net624 vssd1 vssd1 vccd1 vccd1 _02545_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09051__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09239__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10197__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ core.register_file.registers_state\[546\] core.register_file.registers_state\[514\]
+ net688 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08890__B net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _04025_ _04100_ _04203_ _04214_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__o211a_4
XFILLER_0_126_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05322_ _01388_ _01433_ _01434_ _01435_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__or4_1
X_09090_ net2311 net364 net354 _04781_ vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__a22o_1
XANTENNA__06699__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08041_ net485 _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__nor2_1
X_05253_ net1119 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06420__D_N _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05371__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 core.register_file.registers_state\[181\] vssd1 vssd1 vccd1 vccd1 net2221
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 core.register_file.registers_state\[364\] vssd1 vssd1 vccd1 vccd1 net2232
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold924 core.register_file.registers_state\[167\] vssd1 vssd1 vccd1 vccd1 net2243
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11294__RESET_B net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold935 core.register_file.registers_state\[156\] vssd1 vssd1 vccd1 vccd1 net2254
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload36_A clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold946 core.register_file.registers_state\[131\] vssd1 vssd1 vccd1 vccd1 net2265
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06225__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold957 core.register_file.registers_state\[114\] vssd1 vssd1 vccd1 vccd1 net2276
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07422__C1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold968 core.register_file.registers_state\[479\] vssd1 vssd1 vccd1 vccd1 net2287
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ net1479 net540 net519 _02343_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06776__A1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold979 core.register_file.registers_state\[133\] vssd1 vssd1 vccd1 vccd1 net2298
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ net2276 net370 _04935_ net439 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06630__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout299_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ net212 net2332 net371 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
XANTENNA__10005__X _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1006_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _02561_ _03506_ net578 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__o21a_1
XANTENNA__09190__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout466_A _04667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ _03696_ _03860_ _03855_ _03844_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a211o_2
XANTENNA__09478__B1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06707_ net538 _02528_ _02811_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07687_ _01488_ _01550_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__or2_1
XANTENNA__06387__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ net2255 net204 net405 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
X_06638_ net975 _02741_ _02742_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__or3_1
XANTENNA__06161__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__B2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09357_ net1120 net464 _05011_ net415 net1617 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06569_ net968 _02669_ _02672_ _02673_ _02666_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08308_ _01381_ _03140_ net576 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09288_ net1848 _04865_ net337 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
XANTENNA__06805__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09650__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06464__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08239_ _03351_ net575 _04343_ _02488_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10327__S net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11250_ clknet_leaf_68_clk _00762_ net1267 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[722\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ net90 net919 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__and2_1
XANTENNA__06216__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ clknet_leaf_1_clk _00693_ net1137 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[653\]
+ sky130_fd_sc_hd__dfrtp_1
X_10132_ core.pc.current_pc\[28\] _05178_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05975__C1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ net473 _05136_ _05137_ net518 net1550 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06519__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09181__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__C net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08467__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09469__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10965_ clknet_leaf_62_clk _00477_ net1242 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[437\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06378__S0 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08141__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10896_ clknet_leaf_104_clk _00408_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[368\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08991__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06152__C1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11517_ clknet_leaf_18_clk _01029_ net1192 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[989\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08215__B _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold209 core.IO_mod.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11448_ clknet_leaf_3_clk _00960_ net1147 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[920\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09944__A1 core.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ clknet_leaf_11_clk _00891_ net1149 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[851\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05855__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05430__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05940_ core.register_file.registers_state\[302\] core.register_file.registers_state\[270\]
+ core.register_file.registers_state\[430\] core.register_file.registers_state\[398\]
+ net681 net1018 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09172__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1271 net1272 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_68_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1282 net1283 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__clkbuf_4
X_05871_ net954 core.register_file.registers_state\[657\] core.register_file.registers_state\[689\]
+ net709 net646 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a221o_1
XANTENNA__07183__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__B core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07183__B2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1293 net1295 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__clkbuf_4
X_07610_ net449 _03290_ net441 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__or3_1
XANTENNA__10616__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__05590__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ net455 _02717_ net447 vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11090__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08132__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09997__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08683__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ net1052 core.register_file.registers_state\[479\] core.register_file.registers_state\[511\]
+ net679 net1015 vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06143__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09880__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05497__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09211_ net462 net562 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__nand2_4
XFILLER_0_119_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06423_ _01957_ _01987_ _01926_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__or3b_1
XANTENNA__05497__B2 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09227__A3 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09142_ net242 net2409 net349 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__mux2_1
XANTENNA__08435__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06354_ core.register_file.registers_state\[2\] net710 net647 _02458_ vssd1 vssd1
+ vccd1 vccd1 _02459_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_44_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06625__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10242__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05305_ _01405_ _01406_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09073_ net742 net612 net242 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__and3_1
X_06285_ net953 core.register_file.registers_state\[35\] net765 vssd1 vssd1 vccd1
+ vccd1 _02390_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout214_A _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06997__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ _03898_ _04018_ _04126_ _04128_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__a211oi_1
XANTENNA__06997__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold710 core.register_file.registers_state\[438\] vssd1 vssd1 vccd1 vccd1 net2029
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold721 core.register_file.registers_state\[137\] vssd1 vssd1 vccd1 vccd1 net2040
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold732 core.register_file.registers_state\[509\] vssd1 vssd1 vccd1 vccd1 net2051
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08738__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold743 core.register_file.registers_state\[844\] vssd1 vssd1 vccd1 vccd1 net2062
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold754 core.register_file.registers_state\[484\] vssd1 vssd1 vccd1 vccd1 net2073
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 core.register_file.registers_state\[879\] vssd1 vssd1 vccd1 vccd1 net2084
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold776 core.register_file.registers_state\[452\] vssd1 vssd1 vccd1 vccd1 net2095
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold787 core.register_file.registers_state\[892\] vssd1 vssd1 vccd1 vccd1 net2106
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09975_ net1460 core.CPU_DAT_O\[31\] net799 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__mux2_1
Xhold798 core.register_file.registers_state\[453\] vssd1 vssd1 vccd1 vccd1 net2117
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05957__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1231_A core.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05421__A1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ _04785_ net601 vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__nor2_1
XANTENNA__09699__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06299__C net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_X net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09163__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _04889_ net2547 net371 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07174__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08795__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07808_ net514 _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__nor2_1
XANTENNA__08910__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08788_ net565 _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07739_ _03774_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ clknet_leaf_96_clk _00262_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09871__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ net2504 _04889_ net405 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ clknet_leaf_68_clk _00193_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[153\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__A _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold795_A core.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11302_ clknet_leaf_101_clk _00814_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[774\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08729__A2 _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ clknet_leaf_86_clk _00745_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[705\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05946__Y _02051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__B1 _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11164_ clknet_leaf_42_clk _00676_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[636\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ _03945_ _04671_ net556 vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__or3_1
XANTENNA__05412__B2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11095_ clknet_leaf_20_clk _00607_ net1189 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[567\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08986__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05963__A2 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ core.ru.state\[3\] _01443_ _01445_ core.BUSY_O net1129 vssd1 vssd1 vccd1
+ vccd1 _05125_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07165__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06002__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 core.register_file.registers_state\[968\] vssd1 vssd1 vccd1 vccd1 net1389
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 core.register_file.registers_state\[1004\] vssd1 vssd1 vccd1 vccd1 net1400
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08901__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 core.register_file.registers_state\[991\] vssd1 vssd1 vccd1 vccd1 net1411
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_102_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06373__C1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07114__B net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__A1 _04734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ clknet_leaf_80_clk _00460_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[420\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06125__C1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05479__A1 core.decoder.inst\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10879_ clknet_leaf_16_clk _00391_ net1210 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10224__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07130__A _03231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06428__B1 _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06070_ net555 _02147_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__and2_1
XANTENNA__07640__A2 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05651__A1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08599__C _04317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10868__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05585__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout508 net509 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_2
XANTENNA__05403__A1 core.decoder.inst\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06600__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09760_ _04989_ net295 net258 net2043 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06972_ _03075_ _03076_ net970 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__a21o_1
XANTENNA__08896__A _04730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ _04773_ _04774_ _04772_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09145__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05923_ net945 core.register_file.registers_state\[846\] net705 core.register_file.registers_state\[878\]
+ net1018 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a221o_1
X_09691_ net222 net2129 net278 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1090 core.decoder.inst\[16\] vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_33_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08642_ core.IO_mod.data_from_mem\[1\] net246 _04715_ vssd1 vssd1 vccd1 vccd1 _04716_
+ sky130_fd_sc_hd__a21oi_4
X_05854_ net1061 core.register_file.registers_state\[177\] net688 core.register_file.registers_state\[145\]
+ net647 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08573_ net208 _04644_ _04645_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__a31o_1
X_05785_ core.register_file.registers_state\[787\] core.register_file.registers_state\[819\]
+ core.register_file.registers_state\[915\] core.register_file.registers_state\[947\]
+ net695 net652 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__mux4_1
X_07524_ _01613_ _02525_ _03627_ _03628_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__nor4b_1
XTAP_TAPCELL_ROW_46_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08656__A1 core.IO_mod.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07459__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06116__C1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09853__B1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07455_ core.register_file.registers_state\[927\] net700 _03559_ vssd1 vssd1 vccd1
+ vccd1 _03560_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_A _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06406_ net944 core.register_file.registers_state\[449\] net702 core.register_file.registers_state\[481\]
+ net927 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06208__X _02313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07386_ net1108 core.register_file.registers_state\[217\] core.register_file.registers_state\[249\]
+ net858 net829 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ net220 net2399 net349 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__mux2_1
X_06337_ net955 core.register_file.registers_state\[192\] net714 core.register_file.registers_state\[224\]
+ net649 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07092__B1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ net613 net211 vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__and2_1
X_06268_ net952 core.register_file.registers_state\[324\] net710 core.register_file.registers_state\[356\]
+ net1020 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05642__A1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ _03400_ _04110_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold540 core.register_file.registers_state\[620\] vssd1 vssd1 vccd1 vccd1 net1859
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 core.register_file.registers_state\[428\] vssd1 vssd1 vccd1 vccd1 net1870
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06199_ net1049 core.register_file.registers_state\[550\] net750 vssd1 vssd1 vccd1
+ vccd1 _02304_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1126_X net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05495__A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold562 core.register_file.registers_state\[661\] vssd1 vssd1 vccd1 vccd1 net1881
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09384__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 core.register_file.registers_state\[601\] vssd1 vssd1 vccd1 vccd1 net1892
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold584 core.register_file.registers_state\[670\] vssd1 vssd1 vccd1 vccd1 net1903
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 core.register_file.registers_state\[927\] vssd1 vssd1 vccd1 vccd1 net1914
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09958_ core.IO_mod.data_from_mem\[14\] core.CPU_DAT_O\[14\] net800 vssd1 vssd1 vccd1
+ vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XANTENNA__07490__S1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08909_ net573 _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _04982_ net383 net375 net1922 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__a22o_1
XANTENNA__07698__A2 _02630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08895__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07215__A _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ clknet_leaf_28_clk net47 net1195 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10973__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10802_ clknet_leaf_69_clk _00314_ net1273 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[274\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11782_ clknet_leaf_24_clk _01286_ net1183 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08647__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06107__C1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08972__C net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ clknet_leaf_0_clk _00245_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[205\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10664_ clknet_leaf_14_clk _00176_ net1170 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[136\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10595_ clknet_leaf_71_clk _00107_ net1270 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08480__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07622__A2 _03231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11216_ clknet_leaf_104_clk _00728_ net1157 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[688\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09375__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07386__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XANTENNA__07386__B2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
X_11147_ clknet_leaf_109_clk _00659_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[619\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11078_ clknet_leaf_99_clk _00590_ net1166 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[550\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09678__A3 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _01498_ _02560_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__and2_1
XANTENNA__07233__S1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09835__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05570_ _01666_ _01673_ _01674_ _01667_ net932 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_129_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07240_ net808 _03343_ _03344_ net794 vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05872__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05299__B core.decoder.inst\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07171_ net778 _03269_ _03270_ net774 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09063__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06122_ _02219_ _02226_ net1027 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06903__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05624__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06053_ net935 core.register_file.registers_state\[458\] net693 core.register_file.registers_state\[490\]
+ net923 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09366__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06204__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_6
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07916__A3 _02962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09812_ _04711_ _04882_ net458 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__or3b_1
Xfanout327 _05055_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout338 _05046_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_4
Xfanout349 _05025_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_8
X_06955_ core.register_file.registers_state\[554\] core.register_file.registers_state\[522\]
+ net832 vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
X_09743_ _04958_ net290 net275 net1973 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout281_A _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05906_ net951 core.register_file.registers_state\[591\] net709 core.register_file.registers_state\[623\]
+ net660 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a221o_1
XANTENNA__10013__X _05107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _04861_ net287 net282 net2548 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__a22o_1
XANTENNA__10133__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06337__C1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06886_ _02989_ _02990_ net974 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07035__A _03139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ net730 _01489_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nor2_2
X_05837_ net627 _01941_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1190_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06983__S0 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1288_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08556_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__inv_2
X_05768_ net1046 core.register_file.registers_state\[211\] core.register_file.registers_state\[243\]
+ net673 net654 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07507_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__nand2_1
X_08487_ _04562_ _04563_ net600 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07689__B _01550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05699_ net618 _01802_ _01803_ net633 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1076_X net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07438_ _03542_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07369_ net968 _03470_ _03473_ net767 vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_21_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ net2385 net364 net354 _04876_ vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07065__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ net1369 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05615__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09039_ net612 net215 vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__and2_1
XANTENNA__10335__S net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09357__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold370 core.register_file.registers_state\[32\] vssd1 vssd1 vccd1 vccd1 net1689
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold381 net189 vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__B1 core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 core.register_file.registers_state\[659\] vssd1 vssd1 vccd1 vccd1 net1711
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ clknet_leaf_70_clk _00513_ net1275 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[473\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06576__C1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 net852 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06040__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout861 _01458_ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_4
Xfanout872 net874 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_4
Xfanout883 net886 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 _01444_ vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_2
XFILLER_0_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06328__C1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1070 core.register_file.registers_state\[713\] vssd1 vssd1 vccd1 vccd1 net2389
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 core.register_file.registers_state\[594\] vssd1 vssd1 vccd1 vccd1 net2400
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09712__X _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06879__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1092 core.register_file.registers_state\[606\] vssd1 vssd1 vccd1 vccd1 net2411
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11834_ clknet_leaf_36_clk net60 net1224 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09817__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06784__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11765_ clknet_leaf_29_clk _01269_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09293__A1 _04899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11160__RESET_B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10716_ clknet_leaf_40_clk _00228_ net1215 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[188\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11696_ clknet_leaf_70_clk net1508 net1275 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05854__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10647_ clknet_leaf_21_clk _00159_ net1182 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09596__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10578_ clknet_leaf_71_clk _00090_ net1274 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05701__S1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07359__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10363__A0 _05115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05863__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06740_ _02840_ _02844_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09054__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09520__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06671_ net977 _02772_ _02775_ net778 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__a211o_1
XANTENNA__06334__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ net230 _04496_ _04497_ _04500_ _04360_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o32a_1
XFILLER_0_114_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05622_ net1039 core.register_file.registers_state\[727\] core.register_file.registers_state\[759\]
+ net670 net653 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__o221a_1
X_09390_ net1766 net327 net315 _04845_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__a22o_1
XANTENNA__09808__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09070__A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05802__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08341_ _04437_ _04429_ net229 vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05553_ net1039 core.register_file.registers_state\[858\] vssd1 vssd1 vccd1 vccd1
+ _01658_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09284__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06098__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06717__S0 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ core.pc.current_pc\[5\] _04370_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05484_ net1058 core.register_file.registers_state\[348\] vssd1 vssd1 vccd1 vccd1
+ _01589_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07223_ net989 core.register_file.registers_state\[833\] net875 core.register_file.registers_state\[865\]
+ net1075 vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05940__S1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10883__RESET_B net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07047__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11794__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09587__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ _03253_ _03258_ net781 vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06105_ net1046 net751 core.register_file.registers_state\[520\] vssd1 vssd1 vccd1
+ vccd1 _02210_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07085_ net988 core.register_file.registers_state\[70\] net869 core.register_file.registers_state\[102\]
+ net817 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1036_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06270__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06036_ net1036 core.register_file.registers_state\[491\] net747 _02140_ vssd1 vssd1
+ vccd1 vccd1 _02141_ sky130_fd_sc_hd__a31o_1
XANTENNA__09339__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11024__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08011__A2 _04037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06558__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_A net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__X _03422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07987_ _02114_ _03023_ net578 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout663_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06938_ net986 core.register_file.registers_state\[843\] net862 core.register_file.registers_state\[875\]
+ net1069 vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a221o_1
X_09726_ _04924_ net286 net274 net2144 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09511__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A _01459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06869_ net826 _02972_ _02973_ net976 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__o211a_1
X_09657_ _04770_ net286 net282 net1821 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1193_X net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06956__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ net255 _03811_ _04676_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__nor4_1
XANTENNA__08295__S net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09588_ _04941_ net401 net301 net2336 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__a22o_1
XANTENNA__06808__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08539_ core.pc.current_pc\[28\] _04603_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09275__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11550_ clknet_leaf_94_clk _01062_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1022\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07825__A2 _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ clknet_leaf_47_clk _00013_ net1291 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06184__S1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ clknet_leaf_64_clk _00993_ net1249 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[953\]
+ sky130_fd_sc_hd__dfstp_1
Xwire536 _02240_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_4
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09578__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ net1353 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08235__C1 _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ _05115_ net1510 net234 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input57_A gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ net17 net902 net796 net2482 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__o22a_1
XANTENNA__08978__B net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__A0 _02272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06549__C1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07210__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _01514_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout691 net692 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08994__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__A2 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__RESET_B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07403__A _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11817_ clknet_leaf_49_clk _01318_ net1310 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08218__B _03862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09805__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10691__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11748_ clknet_leaf_32_clk _01260_ net1207 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_25_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05827__A1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05827__B2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ clknet_leaf_32_clk _01191_ net1207 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09569__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11047__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09049__B net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__C1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06252__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08888__B net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ net479 _03991_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10336__A0 _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08890_ net226 net739 vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07841_ _03884_ _03916_ _03943_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__and3_1
XANTENNA__07201__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05438__S0 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09065__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06041__X _02146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ core.decoder.inst\[26\] net899 _03875_ _03876_ _03874_ vssd1 vssd1 vccd1
+ vccd1 _03877_ sky130_fd_sc_hd__a221o_2
XANTENNA__05763__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05880__X _01985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ _04771_ net395 net307 net1987 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__a22o_1
X_06723_ core.register_file.registers_state\[786\] core.register_file.registers_state\[818\]
+ core.register_file.registers_state\[914\] core.register_file.registers_state\[946\]
+ net887 net1080 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__mux4_1
XANTENNA__08701__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09442_ _04918_ net315 net311 net1938 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__a22o_1
X_06654_ core.register_file.registers_state\[916\] core.register_file.registers_state\[948\]
+ net888 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11011__RESET_B net1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05605_ net1005 net899 _01507_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ net1762 net329 net321 _04752_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__a22o_1
X_06585_ net552 _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__or2_1
XANTENNA__11831__Q core.IO_mod.input_reg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08324_ core.decoder.inst\[29\] net734 _04420_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_23_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05536_ core.register_file.registers_state\[282\] core.register_file.registers_state\[314\]
+ core.register_file.registers_state\[410\] core.register_file.registers_state\[442\]
+ net696 net1011 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__mux4_1
XANTENNA__08843__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05818__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08255_ _04356_ _04357_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05467_ _01569_ _01571_ net621 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout509_A _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ net994 core.register_file.registers_state\[194\] net884 core.register_file.registers_state\[226\]
+ net815 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06491__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ _03798_ _03879_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__nor2_1
X_05398_ net732 _01496_ _01497_ net724 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08768__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ net815 _03238_ _03237_ net792 vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a211o_1
XANTENNA__06779__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06243__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07068_ _02315_ _02522_ net538 vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout780_A _01462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05451__C1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06019_ core.register_file.registers_state\[811\] core.register_file.registers_state\[779\]
+ net667 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
XANTENNA__10327__A0 _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07194__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__B1 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09709_ net203 net2439 net278 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10981_ clknet_leaf_92_clk _00493_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__C1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11602_ clknet_leaf_24_clk net1619 net1185 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09799__A2 _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07354__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08980__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ clknet_leaf_0_clk _01045_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1005\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06482__A1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05678__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06482__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11464_ clknet_leaf_9_clk _00976_ net1151 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[936\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_115_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07596__C _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08759__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ net1361 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__05690__C1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ clknet_leaf_65_clk _00907_ net1245 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[867\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09420__A1 _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08989__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07893__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10030__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ _05098_ net1521 net232 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07982__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__A0 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ net30 net903 net795 net2528 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__o22a_1
XANTENNA__05993__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09184__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07195__C1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06942__C1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10097__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07498__B1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08229__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09239__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09051__C net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06370_ _02472_ _02473_ net1031 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_100_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05321_ net1122 core.decoder.inst\[8\] core.decoder.inst\[11\] net1116 vssd1 vssd1
+ vccd1 vccd1 _01435_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _03701_ _03723_ net507 vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__mux2_1
XANTENNA__06473__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05252_ net1315 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07670__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06473__B2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold903 core.register_file.registers_state\[837\] vssd1 vssd1 vccd1 vccd1 net2222
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold914 core.register_file.registers_state\[762\] vssd1 vssd1 vccd1 vccd1 net2233
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 core.register_file.registers_state\[503\] vssd1 vssd1 vccd1 vccd1 net2244
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 core.register_file.registers_state\[475\] vssd1 vssd1 vccd1 vccd1 net2255
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08899__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06225__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold947 core.register_file.registers_state\[502\] vssd1 vssd1 vccd1 vccd1 net2266
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 core.register_file.registers_state\[591\] vssd1 vssd1 vccd1 vccd1 net2277
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 core.register_file.registers_state\[340\] vssd1 vssd1 vccd1 vccd1 net2288
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09991_ net1517 net540 net519 net535 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__a22o_1
XANTENNA__10587__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08942_ net571 net216 net738 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__and3_2
XANTENNA__10309__A0 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09175__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09714__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ net205 core.register_file.registers_state\[87\] net371 vssd1 vssd1 vccd1
+ vccd1 _00127_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_68_clk_X clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07824_ core.decoder.inst\[25\] net901 net546 _03928_ vssd1 vssd1 vccd1 vccd1 _03929_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07755_ net511 _03856_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout361_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08135__D1 _02384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_A _05060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06706_ _02526_ _02527_ net538 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__o21a_1
X_07686_ _02518_ _03790_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06387__S1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11212__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ net2479 _04893_ net405 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06637_ net1104 core.register_file.registers_state\[469\] core.register_file.registers_state\[501\]
+ net850 net1077 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ net1115 _05009_ net412 net1902 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a22o_1
X_06568_ net969 _02663_ _02664_ net1066 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__o31a_1
XANTENNA__08426__X _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08307_ core.pc.current_pc\[7\] net598 _04406_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__o21a_1
X_05519_ _01406_ _01490_ _01615_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__or3_1
X_09287_ net2333 net204 net335 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08453__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06499_ _01488_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08238_ core.pc.current_pc\[1\] net575 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__nor2_1
XANTENNA__06464__A1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout995_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05672__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ _01957_ _02900_ net578 vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__o21a_1
XANTENNA__09402__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10200_ net1126 net1613 net911 _05208_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06216__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11180_ clknet_leaf_103_clk _00692_ net1161 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[652\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08602__A _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ _03964_ _05176_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09166__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _04255_ net592 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05727__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__C1 _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10964_ clknet_leaf_55_clk _00476_ net1301 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[436\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06378__S1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ clknet_leaf_84_clk _00407_ net1232 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08991__B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07101__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09641__B2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06455__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ clknet_leaf_44_clk _01028_ net1283 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[988\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_124_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08215__C _04298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11447_ clknet_leaf_8_clk _00959_ net1144 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[919\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06207__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output88_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06731__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ clknet_leaf_64_clk _00890_ net1249 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[850\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07955__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10329_ _05114_ net1740 net239 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05966__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09157__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07128__A _02346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__A1 _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07168__C1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1250 net1278 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_2
Xfanout1261 net1262 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_68_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05870_ core.register_file.registers_state\[529\] core.register_file.registers_state\[561\]
+ net709 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
Xfanout1272 net1277 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__clkbuf_4
Xfanout1283 net1313 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__clkbuf_2
Xfanout1294 net1295 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__clkbuf_2
X_07540_ net552 net443 net451 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__and3b_2
XANTENNA_clkbuf_leaf_80_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09062__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07471_ net1052 core.register_file.registers_state\[351\] core.register_file.registers_state\[383\]
+ net679 net925 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__o221a_1
XANTENNA__09997__B _02204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06143__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08683__A2 _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__B _02145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09880__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06422_ _02016_ _02052_ _02084_ _02114_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__or4_2
XFILLER_0_53_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09210_ _04710_ _04711_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07318__S0 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09141_ net243 net2380 net348 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06353_ net952 core.register_file.registers_state\[34\] net765 vssd1 vssd1 vccd1
+ vccd1 _02458_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_44_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05304_ _01405_ _01406_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__nor2_1
XANTENNA__06446__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ net612 net241 vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__and2_1
XANTENNA__07643__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06284_ core.register_file.registers_state\[163\] net689 net661 _02388_ vssd1 vssd1
+ vccd1 vccd1 _02389_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08023_ net1113 _04125_ _04127_ net578 vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold700 core.register_file.registers_state\[726\] vssd1 vssd1 vccd1 vccd1 net2019
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08199__A1 _03759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout207_A _04705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold711 core.register_file.registers_state\[768\] vssd1 vssd1 vccd1 vccd1 net2030
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__B2 _03771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 core.register_file.registers_state\[224\] vssd1 vssd1 vccd1 vccd1 net2041
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold733 core.register_file.registers_state\[836\] vssd1 vssd1 vccd1 vccd1 net2052
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold744 core.register_file.registers_state\[744\] vssd1 vssd1 vccd1 vccd1 net2063
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 core.register_file.registers_state\[515\] vssd1 vssd1 vccd1 vccd1 net2074
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A1 _02146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 core.register_file.registers_state\[607\] vssd1 vssd1 vccd1 vccd1 net2085
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 core.register_file.registers_state\[252\] vssd1 vssd1 vccd1 vccd1 net2096
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 core.register_file.registers_state\[753\] vssd1 vssd1 vccd1 vccd1 net2107
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ net1453 core.CPU_DAT_O\[30\] net799 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__mux2_1
Xhold799 core.register_file.registers_state\[275\] vssd1 vssd1 vccd1 vccd1 net2118
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1116_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09148__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__S net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__A _03111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ net2457 net368 _04923_ net433 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout576_A _04336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ net741 _04769_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06906__C1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08795__C _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _03910_ _03911_ net488 vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__mux2_1
XANTENNA__05804__S0 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05999_ net617 _02102_ _02103_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout743_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ net605 _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_48_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07738_ _03635_ _03643_ _03708_ _03638_ net479 net490 vssd1 vssd1 vccd1 vccd1 _03843_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__06088__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09320__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout910_A _01449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ net510 _03657_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__nand2_2
XANTENNA__08674__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06134__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__A1 _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09399__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ net2121 _04888_ net406 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06685__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06685__B2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ clknet_leaf_10_clk _00192_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[152\]
+ sky130_fd_sc_hd__dfrtp_1
X_09339_ _04976_ net419 net414 net1663 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a22o_1
XANTENNA__11878__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09623__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07995__X _04100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06117__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout998_X net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ clknet_leaf_101_clk _00813_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[773\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11232_ clknet_leaf_59_clk _00744_ net1286 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[704\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09387__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11163_ clknet_leaf_23_clk _00675_ net1184 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[635\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05948__B1 _01867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09139__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10114_ net1124 core.pc.current_pc\[25\] _05167_ vssd1 vssd1 vccd1 vccd1 _05168_
+ sky130_fd_sc_hd__o21ai_1
X_11094_ clknet_leaf_60_clk _00606_ net1285 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[566\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08986__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ core.ru.state\[0\] _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__nor2_1
XANTENNA__07890__B _03856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold60 core.register_file.registers_state\[1013\] vssd1 vssd1 vccd1 vccd1 net1379
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07382__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 core.register_file.registers_state\[988\] vssd1 vssd1 vccd1 vccd1 net1390
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 core.register_file.registers_state\[1022\] vssd1 vssd1 vccd1 vccd1 net1401
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold93 core.register_file.registers_state\[1008\] vssd1 vssd1 vccd1 vccd1 net1412
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09311__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10947_ clknet_leaf_73_clk _00459_ net1263 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[419\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05479__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07873__B1 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ clknet_leaf_97_clk _00390_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[350\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06428__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__A2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05636__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08242__A _03382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08599__D _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 _02453_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05939__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06061__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05403__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06600__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06971_ net986 core.register_file.registers_state\[458\] net862 core.register_file.registers_state\[490\]
+ net978 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08896__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08710_ core.IO_mod.input_reg\[11\] net253 net727 vssd1 vssd1 vccd1 vccd1 _04774_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__09145__A3 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05922_ net1020 _02026_ _02025_ net934 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a211o_1
X_09690_ _04889_ net2534 net278 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__mux2_1
XANTENNA__06697__A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1080 net1081 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_4
XANTENNA__09550__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__B2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09073__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08641_ core.IO_mod.input_reg\[1\] net250 net725 vssd1 vssd1 vccd1 vccd1 _04715_
+ sky130_fd_sc_hd__a21o_1
X_05853_ net1081 net897 _01867_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10837__RESET_B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06364__B1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08572_ net228 _04646_ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__and3_1
X_05784_ net616 _01887_ _01888_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09302__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07523_ _01550_ _01709_ _02523_ _02533_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_46_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10775__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08656__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07454_ core.register_file.registers_state\[959\] net683 vssd1 vssd1 vccd1 vccd1
+ _03559_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06405_ net944 core.register_file.registers_state\[321\] net702 core.register_file.registers_state\[353\]
+ net1018 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07385_ net1108 core.register_file.registers_state\[89\] core.register_file.registers_state\[121\]
+ net858 net814 vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09605__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09947__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06336_ net956 core.register_file.registers_state\[64\] net715 core.register_file.registers_state\[96\]
+ net663 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a221o_1
X_09124_ _04890_ net2291 net347 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08704__X _04769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09081__A2 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ core.register_file.registers_state\[152\] net427 _05009_ net998 vssd1 vssd1
+ vccd1 vccd1 _00192_ sky130_fd_sc_hd__a22o_1
X_06267_ _02368_ _02371_ net630 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1233_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09369__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08006_ _03400_ _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05642__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06371__S net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 core.register_file.registers_state\[218\] vssd1 vssd1 vccd1 vccd1 net1849
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09908__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08152__A _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06198_ net960 _02297_ _02302_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a21oi_1
Xhold541 core.register_file.registers_state\[770\] vssd1 vssd1 vccd1 vccd1 net1860
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold552 core.register_file.registers_state\[884\] vssd1 vssd1 vccd1 vccd1 net1871
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold563 core.register_file.registers_state\[56\] vssd1 vssd1 vccd1 vccd1 net1882
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 core.register_file.registers_state\[561\] vssd1 vssd1 vccd1 vccd1 net1893
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1021_X net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 core.register_file.registers_state\[51\] vssd1 vssd1 vccd1 vccd1 net1904
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 core.register_file.registers_state\[476\] vssd1 vssd1 vccd1 vccd1 net1915
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1119_X net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__S net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06052__C1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ net1614 core.CPU_DAT_O\[13\] net799 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _04751_ net602 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__nor2_1
X_09888_ _04980_ net386 net378 net1724 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__a22o_1
Xhold1230 net151 vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09541__A0 _04886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ net1121 net604 vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__or2_2
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06355__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08895__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ clknet_leaf_24_clk net45 net1183 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10801_ clknet_leaf_75_clk _00313_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[273\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06107__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout913_X net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ clknet_leaf_29_clk _01285_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08647__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10732_ clknet_leaf_101_clk _00244_ net1163 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[204\]
+ sky130_fd_sc_hd__dfrtp_1
X_10663_ clknet_leaf_91_clk _00175_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[135\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10594_ clknet_leaf_77_clk _00106_ net1262 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07083__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05618__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07885__B _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07083__B2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__05686__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11215_ clknet_leaf_82_clk _00727_ net1232 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[687\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10648__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08997__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06043__C1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09780__B1 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ clknet_leaf_1_clk _00658_ net1133 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[618\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
X_11077_ clknet_leaf_101_clk _00589_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[549\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05625__S net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07406__A _03506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ net1455 net542 net521 _05114_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__a22o_1
XANTENNA__09532__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08099__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07846__A0 _03949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__B2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06456__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06744__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07170_ net1088 _03271_ _03274_ net781 vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05299__C core.decoder.inst\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09063__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06121_ net933 _02220_ _02221_ _02224_ _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__o32a_1
XFILLER_0_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11423__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__RESET_B net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05596__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06052_ net935 core.register_file.registers_state\[330\] net693 core.register_file.registers_state\[362\]
+ net1008 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a221o_1
XANTENNA__06821__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06821__B2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10007__A _01502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 _05064_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09771__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout317 net326 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
X_09811_ net560 _04881_ net461 net272 net1917 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__a32o_1
Xfanout328 _05055_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout339 _05031_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09742_ _04956_ net288 net274 net2263 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a22o_1
X_06954_ core.register_file.registers_state\[618\] core.register_file.registers_state\[586\]
+ net832 vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
XANTENNA__09523__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05905_ _02008_ _02009_ net660 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
XANTENNA__06337__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _04856_ net288 net282 net1934 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__a22o_1
X_06885_ net991 core.register_file.registers_state\[462\] net877 core.register_file.registers_state\[494\]
+ net982 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout274_A _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08624_ net733 _04242_ _01621_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06888__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05836_ _01937_ _01938_ _01939_ _01940_ net1027 net924 vssd1 vssd1 vccd1 vccd1 _01941_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06983__S1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ _04630_ _04631_ _01508_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a21o_1
X_05767_ net1046 core.register_file.registers_state\[83\] core.register_file.registers_state\[115\]
+ net673 net639 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout441_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11877__RESET_B net1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07506_ _03582_ net549 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__nand2_1
X_08486_ _04568_ _04569_ net208 vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05698_ net645 _01790_ _01788_ net618 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05848__C1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07437_ _03511_ _03538_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout706_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1069_X net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11469__SET_B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07368_ net969 _03471_ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_21_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07065__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09107_ net1928 net363 net353 _04871_ vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__a22o_1
X_06319_ net1052 _01408_ _01424_ core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 _02424_
+ sky130_fd_sc_hd__a22oi_4
X_07299_ _02931_ _02934_ _03025_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_111_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1236_X net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06812__A1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09038_ net2370 net430 _04998_ net1000 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06812__B2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold360 core.register_file.registers_state\[918\] vssd1 vssd1 vccd1 vccd1 net1679
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 core.register_file.registers_state\[385\] vssd1 vssd1 vccd1 vccd1 net1690
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06889__X _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 core.register_file.registers_state\[442\] vssd1 vssd1 vccd1 vccd1 net1701
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 core.register_file.registers_state\[411\] vssd1 vssd1 vccd1 vccd1 net1712
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11000_ clknet_leaf_5_clk _00512_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[472\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09762__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10759__RESET_B net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08610__A _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net846 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_2
XANTENNA__10940__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout851 net852 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09109__A3 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout862 net864 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_2
XANTENNA__10351__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 net874 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_2
XANTENNA__08317__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout884 net886 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08317__B2 _04360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05445__S net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09514__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout895 _01410_ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06328__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1060 core.register_file.registers_state\[701\] vssd1 vssd1 vccd1 vccd1 net2379
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 core.register_file.registers_state\[626\] vssd1 vssd1 vccd1 vccd1 net2390
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net1319 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
Xhold1082 core.register_file.registers_state\[148\] vssd1 vssd1 vccd1 vccd1 net2401
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 core.register_file.registers_state\[98\] vssd1 vssd1 vccd1 vccd1 net2412
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07513__X _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__C net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11833_ clknet_leaf_36_clk net57 net1221 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11764_ clknet_leaf_29_clk _01268_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_81_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09293__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10715_ clknet_leaf_19_clk _00227_ net1191 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[187\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_137_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ clknet_leaf_72_clk net1582 net1269 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ clknet_leaf_44_clk _00158_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10577_ clknet_leaf_75_clk _00089_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10060__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06264__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06803__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__B2 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09753__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11129_ clknet_leaf_56_clk _00641_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[601\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09505__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05790__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06670_ _02773_ _02774_ net1089 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__o21a_1
XANTENNA__07531__A2 _02900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05621_ net1039 core.register_file.registers_state\[599\] vssd1 vssd1 vccd1 vccd1
+ _01726_ sky130_fd_sc_hd__or2_1
X_08340_ _04435_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__or2_1
XANTENNA__09070__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05552_ net938 core.register_file.registers_state\[890\] net757 vssd1 vssd1 vccd1
+ vccd1 _01657_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06717__S1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08271_ core.pc.current_pc\[4\] net598 _04373_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05483_ net950 core.register_file.registers_state\[508\] net764 _01587_ net1019 vssd1
+ vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__o311a_1
XFILLER_0_15_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11217__RESET_B net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07222_ net989 core.register_file.registers_state\[961\] net875 core.register_file.registers_state\[993\]
+ net982 vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10813__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07153_ _03254_ _03255_ _03257_ _03256_ net792 net827 vssd1 vssd1 vccd1 vccd1 _03258_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07047__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload59_A clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06104_ net942 core.register_file.registers_state\[552\] net761 vssd1 vssd1 vccd1
+ vccd1 _02209_ sky130_fd_sc_hd__or3_1
XANTENNA__10051__B1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ core.register_file.registers_state\[38\] core.register_file.registers_state\[6\]
+ net842 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06035_ net935 core.register_file.registers_state\[459\] vssd1 vssd1 vccd1 vccd1
+ _02140_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1029_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10852__RESET_B net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout489_A _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ net900 _02085_ net547 _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ _04922_ net289 net275 net1796 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__a22o_1
XANTENNA__11564__Q core.decoder.inst\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06937_ net986 core.register_file.registers_state\[971\] net862 core.register_file.registers_state\[1003\]
+ net978 vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a221o_1
XANTENNA__05781__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _04764_ net291 net283 net2180 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06868_ net1107 core.register_file.registers_state\[686\] core.register_file.registers_state\[654\]
+ net847 net808 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _04028_ _04243_ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__or3_1
XANTENNA__06956__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05819_ _01922_ _01923_ net723 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a21o_1
X_09587_ _04939_ net401 net301 net2258 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout823_A _01459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ _02845_ _02815_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__nand2b_1
X_08538_ net208 _04615_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08469_ _04531_ _04547_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ clknet_leaf_47_clk _00012_ net1291 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05788__X _01893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ clknet_leaf_3_clk _00992_ net1146 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[952\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08605__A _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10431_ net1336 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10346__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10042__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10362_ _05114_ net1759 net235 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10293_ net16 net903 net795 net2436 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__o22a_1
XANTENNA__09735__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08978__C net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 core.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07746__C1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07210__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 net672 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout681 net682 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_4
Xfanout692 _01514_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05772__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05772__B2 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08994__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__A3 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05903__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07390__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__C net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11816_ clknet_leaf_70_clk _01317_ net1276 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11381__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07277__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11747_ clknet_leaf_35_clk _01259_ net1220 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11310__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08074__X _04179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11678_ clknet_leaf_35_clk _01190_ net1220 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10629_ clknet_leaf_87_clk _00141_ net1227 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10033__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06237__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06883__S0 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08888__C net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09726__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08250__A _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07201__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07840_ _03917_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__nor2_1
XANTENNA__05438__S1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06635__S0 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09065__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _01664_ _03476_ net580 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__o21a_1
XANTENNA__05763__A1 core.decoder.inst\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11611__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _04765_ net398 net308 net1925 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__a22o_1
X_06722_ _02823_ _02826_ net774 _02821_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__a211o_2
XANTENNA__08396__S net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _04916_ net319 net312 net2186 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__a22o_1
X_06653_ net828 _02756_ _02757_ net787 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05604_ _01664_ _01708_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09372_ net1992 net328 net318 _04747_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__a22o_1
X_06584_ _01746_ _02688_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09257__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08323_ core.decoder.inst\[29\] net734 _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__and3_1
XANTENNA__07268__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05535_ net621 _01635_ _01636_ _01639_ net628 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_62_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ _04356_ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05466_ core.register_file.registers_state\[29\] net677 net656 _01570_ vssd1 vssd1
+ vccd1 vccd1 _01571_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05401__X _01506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07205_ net994 core.register_file.registers_state\[66\] net884 core.register_file.registers_state\[98\]
+ net830 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a221o_1
X_08185_ _03686_ _04202_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__nor2_1
X_05397_ _01426_ _01489_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__nor2_8
XANTENNA_fanout1146_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07136_ _03239_ _03240_ net787 vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08768__B2 _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11559__Q core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06243__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ net773 _03165_ _03171_ _03160_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__a31o_4
XFILLER_0_112_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1313_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06018_ core.register_file.registers_state\[939\] core.register_file.registers_state\[907\]
+ net667 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XANTENNA__09717__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05784__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10709__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06626__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1101_X net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09690__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__C1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ net530 _04066_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_96_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05754__A1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11291__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09708_ net210 net2355 net281 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
X_10980_ clknet_leaf_75_clk _00492_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09496__A2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__A _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05506__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ _05014_ net396 net391 net2463 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05950__C net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09248__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11601_ clknet_leaf_28_clk _01113_ net1197 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07259__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09799__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07354__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ clknet_leaf_103_clk _01044_ net1155 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1004\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05365__S0 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11463_ clknet_leaf_65_clk _00975_ net1245 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[935\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08759__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__RESET_B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ net1384 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11394_ clknet_leaf_79_clk _00906_ net1253 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[866\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07967__C1 _04070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08989__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07431__A1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10345_ _02272_ net1939 net232 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__mux2_1
XANTENNA__09708__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05442__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08070__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ net29 net904 net797 net2483 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05993__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08931__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05745__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05745__B2 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__A2 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08695__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05320_ net1026 net1053 core.decoder.inst\[24\] vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06317__X _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05356__S0 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__A1_N net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05251_ core.decoder.inst\[14\] vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09947__A0 core.IO_mod.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold904 core.register_file.registers_state\[182\] vssd1 vssd1 vccd1 vccd1 net2223
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold915 core.register_file.registers_state\[574\] vssd1 vssd1 vccd1 vccd1 net2234
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 core.register_file.registers_state\[171\] vssd1 vssd1 vccd1 vccd1 net2245
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08899__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold937 core.register_file.registers_state\[705\] vssd1 vssd1 vccd1 vccd1 net2256
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 core.register_file.registers_state\[201\] vssd1 vssd1 vccd1 vccd1 net2267
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07422__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09990_ net1659 net541 net520 _02421_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__a22o_1
XANTENNA__07422__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold959 core.register_file.registers_state\[662\] vssd1 vssd1 vccd1 vccd1 net2278
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05433__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08941_ net216 net738 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08872_ net741 _04838_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10015__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07186__B1 _01632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07823_ _02561_ _03506_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nand2_1
XANTENNA__08922__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06933__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ net511 _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__nand2_1
XANTENNA__08135__C1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06705_ net771 _02798_ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07489__A1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07685_ net498 _03659_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08686__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10021__Y _05111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout354_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1096_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__RESET_B net1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
X_09424_ net2545 net211 net408 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
X_06636_ net1105 core.register_file.registers_state\[341\] core.register_file.registers_state\[373\]
+ net850 net985 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__o221a_1
XANTENNA__06161__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06161__B2 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ _05007_ net418 net412 net1669 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06567_ net969 _02670_ _02671_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_A _01524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08306_ _04360_ _04405_ _04402_ net209 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05779__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05518_ _01399_ _01614_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__or2_1
XANTENNA__06374__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09286_ net2307 _04893_ net335 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__mux2_1
X_06498_ _01550_ _02602_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__xor2_1
XANTENNA__07110__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09650__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08237_ core.pc.current_pc\[1\] _04335_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__nand2_1
XANTENNA__10260__A3 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05449_ net1043 net749 core.register_file.registers_state\[669\] vssd1 vssd1 vccd1
+ vccd1 _01554_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09938__A0 core.decoder.inst\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09685__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08168_ net901 _01928_ net547 _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout890_A _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout988_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10531__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07119_ net794 _03222_ _03223_ _03221_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a31o_1
X_08099_ _03325_ _03385_ net528 vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a21o_1
XANTENNA__08602__B _04200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10130_ _03964_ _05176_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06621__C1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05975__A1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05975__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__A1 _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10061_ core.pc.current_pc\[4\] net591 vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10681__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__S net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08913__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05727__A1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09469__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11752__Q net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10963_ clknet_leaf_97_clk _00475_ net1168 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[435\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_82_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10894_ clknet_leaf_90_clk _00406_ net1238 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[366\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06152__B2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05360__C1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07101__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09641__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11515_ clknet_leaf_23_clk _01027_ net1184 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[987\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09929__A0 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11446_ clknet_leaf_61_clk _00958_ net1280 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[918\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11377_ clknet_leaf_66_clk _00889_ net1244 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10328_ _05113_ net1519 net239 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
XANTENNA__05966__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05855__C net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10259_ net92 net914 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__and2_1
XANTENNA__07707__A2 _03422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1242 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
Xfanout1251 net1253 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09624__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1262 net1278 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06915__B1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1273 net1277 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__clkbuf_4
Xfanout1284 net1286 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__clkbuf_4
Xfanout1295 net1305 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05590__C net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__C net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_73_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07470_ core.register_file.registers_state\[287\] core.register_file.registers_state\[319\]
+ core.register_file.registers_state\[415\] core.register_file.registers_state\[447\]
+ net700 net1016 vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06143__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07431__X _03536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06421_ _02524_ _02525_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__or2_2
XFILLER_0_118_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09140_ net203 net2428 net348 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__mux2_1
XANTENNA__07318__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06352_ net1059 core.register_file.registers_state\[130\] net688 core.register_file.registers_state\[162\]
+ net661 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__o221a_1
XANTENNA__09093__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05303_ _01417_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ net999 net463 _05019_ net428 net1670 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__a32o_1
X_06283_ net1061 core.register_file.registers_state\[131\] vssd1 vssd1 vccd1 vccd1
+ _02388_ sky130_fd_sc_hd__or2_1
XANTENNA__10242__A3 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08022_ _02241_ _03139_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold701 core.register_file.registers_state\[666\] vssd1 vssd1 vccd1 vccd1 net2020
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold712 core.register_file.registers_state\[213\] vssd1 vssd1 vccd1 vccd1 net2031
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold723 core.register_file.registers_state\[487\] vssd1 vssd1 vccd1 vccd1 net2042
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold734 core.register_file.registers_state\[850\] vssd1 vssd1 vccd1 vccd1 net2053
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 core.register_file.registers_state\[625\] vssd1 vssd1 vccd1 vccd1 net2064
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold756 core.register_file.registers_state\[823\] vssd1 vssd1 vccd1 vccd1 net2075
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold767 core.register_file.registers_state\[741\] vssd1 vssd1 vccd1 vccd1 net2086
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06603__C1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 core.register_file.registers_state\[37\] vssd1 vssd1 vccd1 vccd1 net2097
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ net1548 core.CPU_DAT_O\[29\] net799 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05957__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold789 core.register_file.registers_state\[242\] vssd1 vssd1 vccd1 vccd1 net2108
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05957__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08924_ net568 net206 net736 vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1011_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _04888_ net2112 net372 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout471_A _05127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06906__B1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06877__B net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11413__RESET_B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ _03776_ _03786_ net478 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05804__S1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ net732 _04836_ _04837_ _04835_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a31o_1
XANTENNA__06382__A1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05998_ net1049 core.register_file.registers_state\[204\] core.register_file.registers_state\[236\]
+ net675 net655 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07737_ _02633_ _02634_ _02662_ _03548_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11572__Q core.decoder.inst\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout736_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1099_X net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07668_ net531 _03658_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__nor2_1
XANTENNA__06134__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07341__X _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09871__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09407_ net2188 _04887_ net406 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
X_06619_ core.register_file.registers_state\[533\] core.register_file.registers_state\[565\]
+ net881 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
X_07599_ net502 _03703_ _03702_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05893__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ _04974_ net417 net413 net1665 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a22o_1
XANTENNA__09084__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09623__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ net2081 _04888_ net336 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11300_ clknet_leaf_80_clk _00812_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[772\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06842__C1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08613__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11231_ clknet_leaf_15_clk _00743_ net1214 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[703\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10354__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11162_ clknet_leaf_6_clk _00674_ net1143 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[634\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05948__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08900__X _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ net1124 core.pc.current_pc\[25\] _05092_ vssd1 vssd1 vccd1 vccd1 _05167_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11093_ clknet_leaf_62_clk _00605_ net1242 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[565\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08986__C net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ core.ru.state\[3\] _01445_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_106_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08898__B1 _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold50 core.register_file.registers_state\[10\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold61 core.register_file.registers_state\[989\] vssd1 vssd1 vccd1 vccd1 net1380
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold72 core.register_file.registers_state\[28\] vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 core.register_file.registers_state\[969\] vssd1 vssd1 vccd1 vccd1 net1402
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 core.register_file.registers_state\[1021\] vssd1 vssd1 vccd1 vccd1 net1413
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06373__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05581__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09311__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946_ clknet_leaf_78_clk _00458_ net1252 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[418\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06125__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06125__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05333__C1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ clknet_leaf_18_clk _00389_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[349\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07086__C1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06428__A2 _01745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10224__A3 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_67_clk_X clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ clknet_leaf_100_clk _00941_ net1165 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08050__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05585__C net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__C net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11202__CLK clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ net986 core.register_file.registers_state\[330\] net862 core.register_file.registers_state\[362\]
+ net1069 vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__a221o_1
XANTENNA__06978__A _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07573__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05921_ core.register_file.registers_state\[942\] core.register_file.registers_state\[910\]
+ net687 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08889__B1 _04899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_4
Xfanout1081 core.decoder.inst\[17\] vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08640_ net571 _04707_ net438 net468 net1689 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__a32o_1
X_05852_ net554 _01956_ _01929_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_33_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XANTENNA__09073__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06364__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__A2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ core.pc.current_pc\[30\] _04627_ core.pc.current_pc\[31\] vssd1 vssd1 vccd1
+ vccd1 _04647_ sky130_fd_sc_hd__a21o_1
X_05783_ net1038 core.register_file.registers_state\[851\] core.register_file.registers_state\[883\]
+ net669 net637 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_46_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
X_07522_ _01866_ _02561_ _02598_ _03582_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__or4_1
XANTENNA__06116__A1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06116__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09853__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07453_ net632 _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__nor2_1
X_06404_ net1029 _02508_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07384_ net1108 core.register_file.registers_state\[185\] net858 core.register_file.registers_state\[153\]
+ net813 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a221o_1
XANTENNA__09605__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09123_ net206 net2446 net348 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__mux2_1
X_06335_ _02437_ _02439_ net619 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1059_A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09054_ net742 net462 _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__and3_1
X_06266_ net623 _02369_ _02370_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08005_ _03397_ _03399_ _03142_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_114_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold520 core.register_file.registers_state\[882\] vssd1 vssd1 vccd1 vccd1 net1839
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06197_ net1027 _02299_ _02301_ net933 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a31o_1
Xhold531 core.register_file.registers_state\[38\] vssd1 vssd1 vccd1 vccd1 net1850
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08152__B _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1226_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 core.register_file.registers_state\[548\] vssd1 vssd1 vccd1 vccd1 net1861
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold553 core.register_file.registers_state\[562\] vssd1 vssd1 vccd1 vccd1 net1872
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 core.register_file.registers_state\[870\] vssd1 vssd1 vccd1 vccd1 net1883
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11567__Q core.decoder.inst\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold575 core.register_file.registers_state\[694\] vssd1 vssd1 vccd1 vccd1 net1894
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 core.register_file.registers_state\[524\] vssd1 vssd1 vccd1 vccd1 net1905
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout686_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold597 core.register_file.registers_state\[866\] vssd1 vssd1 vccd1 vccd1 net1916
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09956_ net2092 core.CPU_DAT_O\[12\] net800 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05792__A _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08907_ net2200 net368 _04911_ net433 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__a22o_1
XANTENNA__06240__X _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ _04978_ net386 net375 net1767 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 core.register_file.registers_state\[317\] vssd1 vssd1 vccd1 vccd1 net2539
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1231 core.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07001__C1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ net1847 net467 net434 _04881_ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08769_ core.IO_mod.data_from_mem\[21\] net248 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_101_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ clknet_leaf_104_clk _00312_ net1154 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[272\]
+ sky130_fd_sc_hd__dfrtp_1
X_11780_ clknet_leaf_29_clk _01284_ net1199 vssd1 vssd1 vccd1 vccd1 core.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06107__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08608__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__A3 _04720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07512__A _01399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10731_ clknet_leaf_111_clk _00243_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[203\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10349__S net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05866__B1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10662_ clknet_leaf_96_clk _00174_ net1173 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[134\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10206__A3 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ clknet_leaf_86_clk _00105_ net1228 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__C1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06562__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11225__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10084__S net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11214_ clknet_leaf_82_clk _00726_ net1234 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[686\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08997__B _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06043__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__RESET_B net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
X_11145_ clknet_leaf_38_clk _00657_ net1212 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[617\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07240__C1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__08489__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XANTENNA__07393__S net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__X _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ clknet_leaf_80_clk _00588_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_94_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ net594 _02597_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__nor2_1
XANTENNA__06346__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09296__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09113__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07846__A1 _03950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10929_ clknet_leaf_74_clk _00441_ net1256 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[401\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08237__B _04335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05857__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06120_ net656 _02222_ _02223_ net1007 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_47_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06051_ net958 _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08023__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09220__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10007__B _02051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06034__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ net560 _04877_ net461 net272 net1569 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__a32o_1
Xfanout307 net308 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout318 net320 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout329 _05055_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _04954_ net292 net277 net2026 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06953_ core.register_file.registers_state\[746\] core.register_file.registers_state\[714\]
+ net831 vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__mux2_1
XANTENNA__05793__C1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05904_ core.register_file.registers_state\[687\] core.register_file.registers_state\[655\]
+ net686 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_105_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09672_ _04850_ net297 net284 net2224 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__a22o_1
XANTENNA__10023__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06337__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06884_ net992 core.register_file.registers_state\[334\] net877 core.register_file.registers_state\[366\]
+ net1076 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08623_ core.IO_mod.input_reg\[0\] net249 _04691_ net733 vssd1 vssd1 vccd1 vccd1
+ _04698_ sky130_fd_sc_hd__o211a_1
XANTENNA__09812__A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05835_ net1045 core.register_file.registers_state\[848\] core.register_file.registers_state\[880\]
+ net673 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout267_A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08554_ _01488_ _04335_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10892__CLK clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05766_ net654 _01870_ _01869_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__o21a_1
XANTENNA__08428__A _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _03582_ net549 vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__or2_1
XANTENNA__05404__X _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08485_ _04565_ _04566_ _04567_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11850__Q core.IO_mod.input_reg\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05697_ net659 _01800_ _01801_ _01799_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09958__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1176_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ _03421_ _03422_ _03481_ _03512_ _03540_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08862__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11248__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout601_A _04897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ net1094 core.register_file.registers_state\[602\] core.register_file.registers_state\[634\]
+ net836 net803 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout222_X net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ net2120 net364 net355 _04866_ vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_21_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06318_ net586 _02403_ _02420_ _02387_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_21_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08262__A1 _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07298_ _02999_ _03402_ _03027_ _02937_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ net744 net464 _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06249_ net951 core.register_file.registers_state\[548\] net765 vssd1 vssd1 vccd1
+ vccd1 _02354_ sky130_fd_sc_hd__or3_1
XANTENNA__05615__A3 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1229_X net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09693__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold350 core.register_file.registers_state\[407\] vssd1 vssd1 vccd1 vccd1 net1669
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold361 core.register_file.registers_state\[777\] vssd1 vssd1 vccd1 vccd1 net1680
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold372 core.ru.state\[2\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08565__A2 _01412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__C1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 core.register_file.registers_state\[913\] vssd1 vssd1 vccd1 vccd1 net1702
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold394 core.register_file.registers_state\[796\] vssd1 vssd1 vccd1 vccd1 net1713
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06576__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B1 _03877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 _01459_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
XANTENNA__06576__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout841 net846 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout852 net861 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_2
X_09939_ core.decoder.inst\[28\] core.CPU_DAT_O\[28\] net893 vssd1 vssd1 vccd1 vccd1
+ _01092_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net864 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_4
Xfanout874 _01457_ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_4
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_2
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06328__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1050 core.register_file.registers_state\[338\] vssd1 vssd1 vccd1 vccd1 net2369
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net1318 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
Xhold1061 core.register_file.registers_state\[222\] vssd1 vssd1 vccd1 vccd1 net2380
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 core.register_file.registers_state\[860\] vssd1 vssd1 vccd1 vccd1 net2391
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 core.register_file.registers_state\[180\] vssd1 vssd1 vccd1 vccd1 net2402
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 core.register_file.registers_state\[79\] vssd1 vssd1 vccd1 vccd1 net2413
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11832_ clknet_leaf_28_clk net46 net1194 vssd1 vssd1 vccd1 vccd1 core.IO_mod.input_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11763_ clknet_leaf_37_clk _01267_ net1222 vssd1 vssd1 vccd1 vccd1 core.pc.current_pc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10714_ clknet_leaf_9_clk _00226_ net1152 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[186\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11694_ clknet_leaf_72_clk net1480 net1269 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10645_ clknet_leaf_63_clk _00157_ net1247 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10615__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08073__A _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10576_ clknet_leaf_108_clk _00088_ net1136 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09450__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10060__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06264__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07461__C1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08005__A1 _03397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09202__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08801__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09753__A1 _04975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ clknet_leaf_4_clk _00640_ net1142 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[600\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05775__C1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09505__A1 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06319__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ clknet_leaf_98_clk _00571_ net1169 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[531\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05790__A2 _01893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06319__B2 core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09632__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05620_ net938 core.register_file.registers_state\[631\] net757 vssd1 vssd1 vccd1
+ vccd1 _01725_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09808__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05551_ core.register_file.registers_state\[794\] core.register_file.registers_state\[826\]
+ core.register_file.registers_state\[922\] core.register_file.registers_state\[954\]
+ net696 net1010 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09070__C _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ net230 _04368_ _04369_ _04372_ _04360_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o32a_1
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05482_ net1058 core.register_file.registers_state\[476\] vssd1 vssd1 vccd1 vccd1
+ _01587_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07221_ core.register_file.registers_state\[801\] core.register_file.registers_state\[769\]
+ core.register_file.registers_state\[929\] core.register_file.registers_state\[897\]
+ net849 net1075 vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07152_ core.register_file.registers_state\[932\] core.register_file.registers_state\[900\]
+ net853 vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10051__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06103_ net582 _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05400__A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07083_ net988 core.register_file.registers_state\[166\] core.register_file.registers_state\[134\]
+ net871 net819 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__o221a_1
XANTENNA__09992__B2 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06034_ net935 core.register_file.registers_state\[331\] net1008 vssd1 vssd1 vccd1
+ vccd1 _02139_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06270__A3 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06007__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09744__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06558__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07985_ _02114_ _03023_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout384_A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _04920_ net286 net274 net2191 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__a22o_1
XANTENNA__07688__A1_N core.decoder.inst\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06936_ core.register_file.registers_state\[811\] core.register_file.registers_state\[779\]
+ core.register_file.registers_state\[939\] core.register_file.registers_state\[907\]
+ net832 net1069 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux4_1
XANTENNA__08857__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10821__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _04759_ net290 net282 net2465 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__a22o_1
X_06867_ core.register_file.registers_state\[558\] core.register_file.registers_state\[526\]
+ net847 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08606_ _04064_ _04074_ _04268_ _04680_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05818_ net966 _01919_ net630 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06377__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09586_ _04937_ net397 net302 net1948 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__a22o_1
X_06798_ _02875_ _02902_ _02876_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__o21a_1
XANTENNA__06191__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08537_ _04607_ _04614_ _04613_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a21o_1
XANTENNA__11070__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11580__Q core.decoder.inst\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05749_ net1064 core.register_file.registers_state\[340\] core.register_file.registers_state\[372\]
+ net691 net929 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1081_X net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_X net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09688__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07997__A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10638__CLK clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _01747_ _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__xor2_1
XANTENNA__09680__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06494__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07419_ net1091 core.register_file.registers_state\[184\] net831 core.register_file.registers_state\[152\]
+ net802 vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08399_ core.pc.current_pc\[16\] net577 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire549 _03606_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__buf_4
X_10430_ net1323 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08235__A1 _03319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05310__A core.control_logic.instruction\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ _05113_ net1562 net235 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__mux2_1
XANTENNA__10042__B2 _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07936__S net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08180__X _04285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ net15 net904 _05244_ core.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 _01289_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08621__A _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10362__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 core.CPU_DAT_I\[28\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 net156 vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06549__A1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 net663 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout671 net672 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout682 net685 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_8
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08710__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06182__C1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11815_ clknet_leaf_70_clk _01316_ net1274 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10110__B net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11768__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11746_ clknet_leaf_35_clk _01258_ net1220 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09671__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10281__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06485__B1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11677_ clknet_leaf_35_clk _01189_ net1220 vssd1 vssd1 vccd1 vccd1 core.ADR_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ clknet_leaf_75_clk _00140_ net1259 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06316__A _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10033__A1 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10559_ clknet_leaf_94_clk _00071_ net1176 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06883__S1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06051__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__S0 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06635__S1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ net1114 _03873_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__or2_1
XANTENNA__05763__A2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06986__A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06721_ net977 _02824_ _02825_ net782 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__o31a_1
XANTENNA__11093__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08701__A2 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _04914_ net320 net312 net2325 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__a22o_1
X_06652_ net996 core.register_file.registers_state\[660\] core.register_file.registers_state\[692\]
+ net889 net814 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a221o_1
X_05603_ net555 _01688_ _01706_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__o31a_2
XFILLER_0_93_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09371_ net2207 net328 net318 _04742_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__a22o_1
X_06583_ net539 _01781_ _02687_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a21o_1
X_08322_ core.pc.current_pc\[9\] _03111_ net576 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05534_ net653 _01637_ _01638_ net616 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_62_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09662__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload71_A clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06476__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ _04340_ _04350_ _04339_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a21o_1
X_05465_ net1051 core.register_file.registers_state\[61\] net751 vssd1 vssd1 vccd1
+ vccd1 _01570_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10930__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07204_ _03306_ _03308_ net787 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08184_ _02906_ _03410_ _02847_ _02903_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05396_ _01399_ _01496_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nand2_1
XANTENNA__10019__Y _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06228__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09965__A1 core.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__B2 _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07135_ net994 core.register_file.registers_state\[196\] net884 core.register_file.registers_state\[228\]
+ net815 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__a221o_1
XANTENNA__08768__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1041_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06779__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06779__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07066_ net1086 _03169_ _03170_ net1067 _03168_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a311o_1
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05987__C1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05451__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05451__B2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06017_ _02118_ _02119_ _02120_ _02121_ net620 net651 vssd1 vssd1 vccd1 vccd1 _02122_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10035__X _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1306_A net1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09971__S net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05739__C1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06626__S1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11436__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A _01509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08940__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _03657_ _03860_ _04072_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_138_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06919_ _02114_ _02932_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__xor2_1
X_09707_ net204 net2552 net278 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
X_07899_ net529 _03988_ _03989_ _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout933_A _01375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1296_X net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _05013_ net396 net392 net2020 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06703__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06164__C1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _04903_ net402 net300 net2158 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11600_ clknet_leaf_28_clk _01112_ net1198 vssd1 vssd1 vccd1 vccd1 core.IO_mod.data_from_mem\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08175__X _04280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09653__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ clknet_leaf_110_clk _01043_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[1003\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_37_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06467__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__S net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05365__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11462_ clknet_leaf_99_clk _00974_ net1159 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[934\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09956__A1 core.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__A2 _04317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ net1328 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__05690__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11393_ clknet_leaf_86_clk _00905_ net1225 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[865\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07967__B1 _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input62_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ _02314_ net1559 net234 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05442__A1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10275_ net28 net903 net795 core.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_128_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09184__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__B2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08931__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06942__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06942__B2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10953__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08447__A1 _04515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09644__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09121__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10254__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11729_ clknet_leaf_45_clk _01241_ net1288 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05356__S1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05250_ net1114 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkinv_4
XANTENNA__07670__A2 _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05681__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09947__A1 core.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10006__B2 _05103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold905 core.register_file.registers_state\[697\] vssd1 vssd1 vccd1 vccd1 net2224
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold916 core.register_file.registers_state\[799\] vssd1 vssd1 vccd1 vccd1 net2235
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 core.register_file.registers_state\[709\] vssd1 vssd1 vccd1 vccd1 net2246
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 core.register_file.registers_state\[332\] vssd1 vssd1 vccd1 vccd1 net2257
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05969__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold949 core.register_file.registers_state\[846\] vssd1 vssd1 vccd1 vccd1 net2268
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11459__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ net2383 net370 _04933_ net438 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09175__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08871_ _04832_ net2001 net373 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10015__B _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07186__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07822_ net489 _03926_ _03924_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_4_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08922__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10190__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06933__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _03720_ _03825_ _03857_ net489 vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ net780 _02803_ _02808_ net767 vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__o211a_1
X_07684_ _01488_ net450 net442 net505 vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__o31a_1
XANTENNA__10031__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09883__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ net2381 net212 net405 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
XANTENNA__11531__SET_B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06635_ core.register_file.registers_state\[277\] core.register_file.registers_state\[309\]
+ core.register_file.registers_state\[405\] core.register_file.registers_state\[437\]
+ net881 net1077 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout347_A _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1089_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ net1120 _05006_ net415 net1616 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__a22o_1
XANTENNA__06655__S net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06566_ net1094 core.register_file.registers_state\[599\] core.register_file.registers_state\[631\]
+ net835 net803 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08305_ _04403_ _04404_ net598 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__o21a_1
X_05517_ core.decoder.inst\[30\] _01618_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09285_ net2405 net211 net338 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__mux2_1
X_06497_ _01613_ net537 _02601_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07110__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout514_A _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1256_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ _04339_ _04340_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09966__S net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05448_ net942 core.register_file.registers_state\[573\] net761 vssd1 vssd1 vccd1
+ vccd1 _01553_ sky130_fd_sc_hd__or3_1
XANTENNA__08723__X _04785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05672__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08167_ _01957_ _02900_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05379_ core.register_file.registers_state\[542\] core.register_file.registers_state\[574\]
+ net876 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_X net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07118_ net990 core.register_file.registers_state\[197\] net876 core.register_file.registers_state\[229\]
+ net809 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08098_ _04017_ _04202_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout883_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08602__C _04215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__A3 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07049_ net794 _03152_ _03153_ net783 vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10826__CLK clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ net473 _05134_ _05135_ net517 net1599 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__A2 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06385__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08677__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ clknet_leaf_69_clk _00474_ net1266 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[434\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09874__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10893_ clknet_leaf_0_clk _00405_ net1132 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[365\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06783__S0 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06418__X _02523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10236__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07101__A1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11514_ clknet_leaf_6_clk _01026_ net1145 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[986\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_136_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11445_ clknet_leaf_63_clk _00957_ net1241 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[917\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10995__RESET_B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07396__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11376_ clknet_leaf_105_clk _00888_ net1156 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[848\]
+ sky130_fd_sc_hd__dfrtp_1
X_10327_ _05112_ net1475 net240 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09157__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ net1125 net1484 net910 _05237_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__a31o_1
XANTENNA__07168__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1230 net1232 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08904__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
X_10189_ net117 net919 net908 net1455 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a22o_1
Xfanout1252 net1253 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10172__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1263 net1268 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1274 net1276 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09116__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1285 net1286 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__clkbuf_4
Xfanout1296 net1305 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08668__B2 _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09865__B1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__X _03817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09640__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__A3 _03763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07340__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06420_ _02146_ _02206_ _02241_ _02176_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__or4b_1
XANTENNA__09880__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09617__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06351_ net554 _02455_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05302_ _01408_ net895 _01416_ _01397_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__and4b_2
XTAP_TAPCELL_ROW_44_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09070_ net746 net612 _04875_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06282_ net586 _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07643__A2 _03052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08021_ net546 _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11281__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05654__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08703__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold702 core.register_file.registers_state\[437\] vssd1 vssd1 vccd1 vccd1 net2021
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 core.register_file.registers_state\[876\] vssd1 vssd1 vccd1 vccd1 net2032
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09396__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold724 core.register_file.registers_state\[782\] vssd1 vssd1 vccd1 vccd1 net2043
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold735 core.register_file.registers_state\[518\] vssd1 vssd1 vccd1 vccd1 net2054
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload34_A clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold746 core.register_file.registers_state\[564\] vssd1 vssd1 vccd1 vccd1 net2065
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold757 core.register_file.registers_state\[686\] vssd1 vssd1 vccd1 vccd1 net2076
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold768 core.register_file.registers_state\[318\] vssd1 vssd1 vccd1 vccd1 net2087
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ net1611 core.CPU_DAT_O\[28\] net799 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__mux2_1
Xhold779 core.register_file.registers_state\[232\] vssd1 vssd1 vccd1 vccd1 net2098
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09148__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ _04780_ net736 vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__and2_1
XANTENNA__10999__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net741 _04763_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1004_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06367__C1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ _03784_ _03801_ net481 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11853__Q core.IO_mod.input_reg\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08785_ core.IO_mod.data_from_mem\[23\] net247 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nand2_1
X_05997_ net1049 core.register_file.registers_state\[76\] core.register_file.registers_state\[108\]
+ net675 net640 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__o221a_1
XFILLER_0_137_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06382__A2 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ _02662_ _03548_ _02633_ _02634_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06119__C1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09856__B1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _03759_ _03771_ net510 vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout631_A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ net1885 _04886_ net407 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__mux2_1
X_06618_ _02721_ _02722_ net794 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07882__A2 _03412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ net454 _03111_ net446 vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__and3_1
XANTENNA__08166__A _03685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06238__X _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10218__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07070__A _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09337_ _04972_ net419 net412 net1643 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__a22o_1
X_06549_ net810 _02652_ _02653_ net1087 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a211o_1
XANTENNA__11624__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09696__S net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05302__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ net2321 _04887_ net336 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ net255 _03811_ _04322_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__nand4_1
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06117__C net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07871__A2_N net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06842__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09199_ _05003_ net358 net425 net1824 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__a22o_1
XANTENNA__08613__B _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ clknet_leaf_96_clk _00742_ net1178 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09387__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06414__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ clknet_leaf_56_clk _00673_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[633\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05948__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10112_ net470 _05165_ _05166_ net515 net1437 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11092_ clknet_leaf_56_clk _00604_ net1293 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[564\]
+ sky130_fd_sc_hd__dfrtp_1
X_10043_ _01438_ net556 core.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__and3b_1
XANTENNA__07516__Y _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 core.register_file.registers_state\[997\] vssd1 vssd1 vccd1 vccd1 net1359
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold51 core.register_file.registers_state\[1002\] vssd1 vssd1 vccd1 vccd1 net1370
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold62 core.register_file.registers_state\[975\] vssd1 vssd1 vccd1 vccd1 net1381
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 core.register_file.registers_state\[24\] vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 core.register_file.registers_state\[986\] vssd1 vssd1 vccd1 vccd1 net1403
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 core.register_file.registers_state\[973\] vssd1 vssd1 vccd1 vccd1 net1414
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_19_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11154__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__B1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09311__A2 _04933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10945_ clknet_leaf_83_clk _00457_ net1230 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11123__RESET_B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__A2_N net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07873__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ clknet_leaf_43_clk _00388_ net1282 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[348\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07086__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08804__A core.IO_mod.input_reg\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05636__B2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09378__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11428_ clknet_leaf_80_clk _00940_ net1254 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[900\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11359_ clknet_leaf_15_clk _00871_ net1177 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[831\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09635__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05920_ _02023_ _02024_ net929 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08889__B2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05851_ _01936_ _01942_ _01949_ _01955_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__o22a_4
XANTENNA_clkbuf_leaf_6_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1083 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1093 net1103 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_4
X_08570_ core.pc.current_pc\[30\] core.pc.current_pc\[31\] _04627_ vssd1 vssd1 vccd1
+ vccd1 _04646_ sky130_fd_sc_hd__nand3_1
X_05782_ net1038 core.register_file.registers_state\[979\] core.register_file.registers_state\[1011\]
+ net669 net652 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__o221a_1
XANTENNA__09838__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ _02604_ _03550_ _03614_ net527 vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09302__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11647__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07452_ _03553_ _03554_ _03555_ _03556_ net622 net642 vssd1 vssd1 vccd1 vccd1 _03557_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06521__C1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06403_ core.register_file.registers_state\[289\] core.register_file.registers_state\[257\]
+ core.register_file.registers_state\[417\] core.register_file.registers_state\[385\]
+ net681 net1017 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07383_ net829 _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09066__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09122_ net222 net2544 net347 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
X_06334_ core.register_file.registers_state\[0\] net714 net649 _02438_ vssd1 vssd1
+ vccd1 vccd1 _02439_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06824__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09053_ net612 _04844_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06265_ net953 core.register_file.registers_state\[196\] net710 core.register_file.registers_state\[228\]
+ net647 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout212_A _04844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ net529 _04045_ _04097_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a31o_2
XFILLER_0_103_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09369__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold510 core.register_file.registers_state\[767\] vssd1 vssd1 vccd1 vccd1 net1829
+ sky130_fd_sc_hd__dlygate4sd3_1
X_06196_ net1045 core.register_file.registers_state\[998\] net750 _02300_ net924 vssd1
+ vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a311o_1
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 core.register_file.registers_state\[789\] vssd1 vssd1 vccd1 vccd1 net1840
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 core.register_file.registers_state\[559\] vssd1 vssd1 vccd1 vccd1 net1851
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 core.register_file.registers_state\[899\] vssd1 vssd1 vccd1 vccd1 net1862
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 core.register_file.registers_state\[566\] vssd1 vssd1 vccd1 vccd1 net1873
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 core.register_file.registers_state\[237\] vssd1 vssd1 vccd1 vccd1 net1884
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__C1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1121_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 core.register_file.registers_state\[751\] vssd1 vssd1 vccd1 vccd1 net1895
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1219_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 core.register_file.registers_state\[853\] vssd1 vssd1 vccd1 vccd1 net1906
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 core.register_file.registers_state\[831\] vssd1 vssd1 vccd1 vccd1 net1917
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ net1594 core.CPU_DAT_O\[11\] net800 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net568 _04746_ net736 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and3_1
XANTENNA__10136__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _04976_ net387 net376 net2136 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__a22o_1
Xhold1210 core.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1007_X net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1221 core.register_file.registers_state\[96\] vssd1 vssd1 vccd1 vccd1 net2540
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 core.pc.current_pc\[13\] vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11583__Q core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ net568 net607 net242 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__and3_1
XANTENNA__10203__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_A _01458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__A0 _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ net2006 net469 net439 _04822_ vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__a22o_1
X_07719_ net482 _03821_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08699_ net567 _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__and2_1
XANTENNA__08608__B _03811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ clknet_leaf_111_clk _00242_ net1131 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[202\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ clknet_leaf_100_clk _00173_ net1164 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07068__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10592_ clknet_leaf_52_clk _00104_ net1303 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05618__B2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10365__S net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11213_ clknet_leaf_2_clk _00725_ net1148 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_92_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08032__A2 _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06579__C1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08630__Y _04705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06043__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ clknet_leaf_13_clk _00656_ net1171 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[616\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09780__A2 _04707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ clknet_leaf_66_clk _00587_ net1264 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[547\]
+ sky130_fd_sc_hd__dfrtp_1
X_10026_ net1488 net542 net521 _05113_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__a22o_1
XANTENNA__09532__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__CLK clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__RESET_B net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06751__C1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09296__A1 _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10928_ clknet_leaf_108_clk _00440_ net1140 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[400\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06503__C1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10859_ clknet_leaf_110_clk _00371_ net1130 vssd1 vssd1 vccd1 vccd1 core.register_file.registers_state\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07059__B1 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05609__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08271__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06050_ core.register_file.registers_state\[298\] core.register_file.registers_state\[266\]
+ core.register_file.registers_state\[426\] core.register_file.registers_state\[394\]
+ net669 net1009 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_10_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10366__A0 _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06989__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09365__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 _05063_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_4
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07156__Y _03261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ _04952_ net287 net274 net2373 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__a22o_1
X_06952_ core.register_file.registers_state\[682\] core.register_file.registers_state\[650\]
+ net834 vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
.ends

